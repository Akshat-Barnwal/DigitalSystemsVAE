`timescale 1s/1ps
module layer6(clk,reset,x,y,done);
input clk,reset;
output done;
input signed [17:0]x[0:19];
output signed [17:0]y[0:783];
localparam signed [17:0]W[0:15679] = {
-24506,-15490,-15491,-5443,-13291,-20799,-3050,-22692,-11302,-7122,-20155,-23644,-7106,-6224,-19761,-16366,-38159,-14262,-29256,-6904,
-27894,-7974,-23581,-10091,-11258,-19925,-8045,-30910,-3629,-10324,-17344,-26118,-15320,-9090,-21762,-14266,-41437,-12711,-22612,-14410,
-23095,-9300,-19179,-6853,-13738,-18071,-6964,-19955,-4013,-15289,-19306,-17305,-18764,-7354,-21628,-10341,-38606,-16043,-27117,-9647,
-18496,-9004,-15633,-13809,-20570,-24982,-13037,-27635,-12553,-15098,-17703,-21316,-17992,-3311,-10377,-8562,-33730,-20233,-20192,-5442,
-24451,-9257,-23147,-13183,-10549,-21275,-6972,-38127,-13674,-15444,-23611,-35908,-14647,-7263,-16155,-14637,-36525,-15549,-16650,-9144,
-21839,-14968,-13080,-9501,-12040,-25695,-8302,-19024,-11719,-15251,-15228,-18117,-5081,-4371,-18882,-4349,-37596,-13540,-34994,-11892,
-24772,-5672,-11459,-16205,-15868,-32616,-12973,-15011,-10017,-7930,-11333,-10175,-9385,-5736,-18800,-3716,-38117,-7026,-29530,-11114,
-23693,-4640,-12299,-7983,-21497,-21450,-3029,-15555,-2958,-10294,-8372,-17042,-15286,-8837,-20352,-14925,-43489,-4971,-27140,-5079,
-20608,-16001,-21019,-8927,-21715,-17257,-7906,-22416,-3347,-8781,-6493,-20473,-11382,-5643,-23788,-2760,-40323,-17752,-32496,-13182,
-23938,-4173,-13161,-6120,-18138,-20682,-9349,-22644,-7201,-16761,-18543,-16056,-6298,-7421,-21687,-14502,-39326,-12399,-28007,-7947,
-24516,-13657,-13942,-4288,-13438,-19577,-8056,-19267,-15033,-20196,-10790,-18090,-6117,-5642,-19644,-10751,-37160,-5901,-33163,-7954,
-19343,-5582,-19659,-7093,-17322,-19120,-376,-14765,-3106,-8916,-11875,-25775,-16570,-8381,-21059,-15373,-39032,-15628,-22421,-13302,
-22785,-5396,-20288,-11558,-19433,-15508,-2815,-31260,-6745,-19053,-21480,-17483,-15658,-11176,-18913,-10340,-28437,-12950,-28386,-16605,
-28341,-16757,-12361,-14212,-13154,-13966,-10995,-20545,-13120,-17371,-27996,-33308,-7441,-16905,-13905,-17323,-28878,-6135,-19654,-7792,
-21179,-4839,-8563,-11297,-22070,-10470,-9205,-24988,-15506,-20017,-21992,-31210,-7853,-15278,-12402,-10534,-27236,-11207,-26449,-11730,
-29169,-12647,-10466,-6262,-13578,-20113,-3287,-30287,-7583,-12076,-18401,-18477,-15059,-12841,-22824,-12746,-37739,-19499,-23529,-7697,
-17394,-10784,-15702,-10697,-17658,-24435,-4449,-21688,-6972,-13654,-12202,-19399,-11590,-10990,-23582,-7155,-44297,-6285,-24966,-10616,
-16520,-3452,-19851,-12447,-19825,-28355,-8262,-12885,-3423,-8950,-6746,-17798,-12052,-3400,-19483,-11431,-42505,-5035,-29983,-11075,
-14571,-11746,-20925,-5994,-16596,-28951,-5588,-23970,-11324,-17530,-11350,-16845,-10859,-4823,-16903,-9843,-36207,-5074,-26779,-17436,
-29490,-12034,-13828,-13527,-10161,-14275,-13224,-39017,-13262,-22004,-16713,-38850,-16899,-11392,-9849,-15825,-34984,-13882,-20901,-20480,
-23597,-3777,-9076,-2278,-18835,-24046,-7876,-18385,-7897,-5836,-17760,-19028,-7056,-10420,-16459,-15481,-34447,-8727,-30338,-5684,
-17748,-7875,-9979,-13511,-11936,-24030,-10354,-40081,-14493,-23211,-12349,-22342,-15208,-6993,-13657,-11777,-39491,-14724,-27253,-11200,
-20172,-7332,-16357,-15950,-21005,-26071,-13039,-16990,-6811,-12367,-9265,-27020,-7530,-13932,-18789,-2672,-39145,-11725,-28207,-12916,
-21173,-9703,-18872,-13032,-21277,-26044,-8673,-23171,-4143,-11106,-10998,-22886,-11283,-13018,-21980,-2512,-36020,-13108,-31625,-11905,
-25953,-10565,-12160,-7936,-13424,-18161,-6232,-26832,-13775,-11738,-21904,-24322,-13380,-18801,-10053,-16183,-35497,-19827,-27579,-10231,
-20715,-10205,-15468,-5474,-16238,-22833,-974,-12428,-6314,-13784,-16181,-11190,-9597,-15682,-25915,-4021,-40925,-5876,-34472,-12546,
-16732,-6606,-18768,-8481,-18357,-23328,214,-23031,-3285,-10660,-16145,-9200,-14688,-8617,-25111,-12853,-34963,-5066,-35228,-5463,
-22265,-4535,-14167,-9388,-19523,-17618,-12706,-37029,-14464,-23253,-14203,-25328,-16301,-15085,-15284,-4140,-31706,-11302,-30115,-10972,
-13670,-8049,-13978,-4539,-18899,-24612,-5755,-14397,-6012,-10190,-6114,-15169,-12761,-6033,-26083,-10660,-46389,-5573,-29908,-8387,
-25617,-16774,-10283,-13748,-15628,-22613,-4153,-19179,-8803,-8739,-18401,-17181,-6375,-18085,-20987,-13993,-44772,-15002,-24939,-7716,
-21203,-2550,-14604,-4231,-20331,-19764,-5668,-12429,-7161,-6700,-16915,-22100,-4895,-8610,-21092,-12691,-41930,-15077,-29677,-2788,
-15477,-1981,-18961,-5546,-15944,-26620,-239,-17425,-6980,-7872,-7918,-20956,-9385,-8631,-26043,-5773,-42179,-5799,-33440,-2010,
-21021,-9152,-13512,-9859,-16226,-18338,-1946,-29790,-11894,-21192,-17869,-20728,-19067,-6444,-16969,-8106,-36924,-13428,-25248,-6413,
-19203,-3160,-13859,-14050,-12344,-27338,-11458,-20519,-7054,-12419,-16901,-16239,-14164,-6827,-21693,-4781,-32582,-15958,-28102,-12634,
-20028,-5954,-8287,-17451,-7481,-22371,-9715,-32624,-5887,-23085,-16964,-19710,-13136,-12655,-17557,-15124,-30207,-15981,-19192,-8099,
-12427,-2277,-16273,-8974,-14258,-17923,-4870,-24801,-5642,-11616,-1247,-20924,-8864,-15899,-25753,-15124,-29421,-10171,-16587,-11206,
-11145,-13826,-13688,-15179,-17581,-9766,-9540,-28568,-11191,-14074,2250,-20850,-6514,-11508,-22432,-10250,-21681,-17269,-13188,-10018,
-12272,-17891,-19167,-15058,-8132,-9260,-11477,-22697,-21746,-15220,-907,-18057,-16579,-13000,-21482,-5113,-18605,-14997,-8907,-7820,
-15011,-16456,-14362,-14088,-16611,-9925,-13897,-8154,-10351,-12124,4145,-12875,-7179,-12022,-27499,-6966,-11471,-7120,-19464,-15193,
-19713,-15723,-10213,-17498,-7027,-19368,-5263,-6560,-14818,-9828,-590,-20795,-3562,-8247,-22993,-5280,-9398,-4028,-21697,-5112,
-37853,-9269,-15495,-16927,-17826,-15745,-12230,-11682,-20923,-7535,-7997,-12431,-7814,-1658,-24030,-4542,-9594,-5120,-10381,-782,
-40626,-23167,-13954,-5928,-8188,-15740,-10571,-9464,-29929,164,-24357,-9631,-13740,2193,-14586,-16331,-5214,-9847,-15993,1553,
-47151,-18978,-1008,-10682,-20794,-15612,-15861,-9157,-20847,-1324,-26707,-19260,-16715,-2823,-20573,-15751,-3314,-5675,-15424,-1428,
-60221,-16401,-12787,-13097,-21252,-17139,-4568,-5805,-11110,4195,-17316,-7441,-12536,-8933,-25866,-12170,-3967,344,-23458,2033,
-50512,-10908,-9107,-13249,-23707,-23836,-8009,-1384,-22926,3765,-28550,-8928,-9913,-9162,-17920,-11565,-7384,-9310,-11969,8218,
-43231,-18099,-15307,-11957,-14640,-18505,-8627,-2006,-29235,8232,-34760,-8295,-16997,251,-12605,-10594,-5531,-10288,-22393,7889,
-42261,-11349,-5522,-5172,-30899,-22617,-15453,3773,-14193,-130,-22468,-22912,-7015,-4398,-19394,-9633,-8868,-6614,-24112,2673,
-34496,4301,-3900,-12529,-24124,-21047,-4962,-2297,-21405,-1945,-50742,-16759,-10249,-3677,-15779,-18194,-13312,-4576,-19276,5252,
-35350,-4236,-6130,-5633,-25080,-26347,-9238,-7788,-18313,6599,-51673,-23522,-12127,-7601,-19638,-7916,-8698,-5231,-22451,4325,
-34104,-6998,-11293,-11253,-17812,-24558,-7307,-14855,-6362,-7073,-17507,-15467,-13292,-5027,-25250,-5765,-12035,-11561,-27322,4040,
-24534,-5096,-6064,-8664,-23781,-21188,-5912,-11050,-5553,-3516,-13094,-21950,-13855,-8568,-17083,-14099,-27057,-3368,-24360,-4329,
-25858,-10319,-20603,-4183,-18794,-27026,-5919,-31079,-6262,-19525,-22621,-18895,-4725,-16645,-26333,-5398,-31614,-16960,-21227,-14158,
-22197,-4214,-11728,-5750,-13890,-19989,-1857,-19736,-13394,-17606,-13288,-15579,-7650,-4660,-19620,-15923,-37096,-15447,-32800,-17826,
-26517,-14415,-21988,-8978,-20004,-12240,-8577,-34407,-16265,-18403,-20009,-21386,-11626,-5468,-11730,-13753,-37882,-17278,-19974,-6413,
-17880,-12091,-9839,-9072,-13288,-28150,-897,-25472,-15206,-7799,-19572,-15685,-16238,-6026,-13760,-5422,-34275,-4483,-31212,-12848,
-25907,-14304,-14349,-6192,-13250,-16796,-6883,-31664,-4757,-20047,-16919,-30678,-18934,-6201,-21242,-11671,-32726,-16592,-29243,-7557,
-22797,-9581,-17124,-7940,-22596,-21918,-10033,-10376,-7792,-5746,-14953,-14399,-10651,-4501,-17157,-8124,-35167,-13050,-32822,-2953,
-17088,-1252,-13961,-4665,-13868,-20626,-2053,-15607,-9208,-16398,-5901,-23981,-5362,-8335,-24466,-7276,-44144,-12978,-36400,-7865,
-23546,-13320,-11841,-5807,-23009,-24044,-51,-20855,-8552,-15613,-14856,-22807,-4215,-7536,-19000,-11447,-28010,-18185,-31389,-14230,
-26592,-2117,-19982,-12313,-18819,-23468,-7088,-25609,-3027,-8235,-9624,-23007,-9469,-8437,-19399,-5198,-31476,-17193,-28174,-9507,
-25134,-4585,-13917,-4114,-18776,-22067,-10370,-10534,-9342,-3795,-20572,-26070,-12277,-10956,-18223,-12273,-27276,-15203,-18566,-2209,
-23629,-4303,-16185,-15167,-12061,-25432,-11513,-16416,-5407,-8814,-8161,-15433,-13191,-15721,-22425,-3588,-33544,-10229,-26910,-4261,
258,-7261,-13952,-10249,-8346,-16981,-540,-11194,-15410,-8520,1695,-17112,-11753,-3631,-22413,-6356,-19693,-15822,-17865,-6278,
-1765,-3533,-13922,-10035,-7994,-8114,-10544,-25613,-17321,-15571,-6015,-12759,-16385,-12096,-26474,-6200,-9661,-4494,-18536,-11554,
-3483,-18274,-4563,-18342,-5988,-12034,-3060,-23784,-23404,-6985,-3837,-19550,-4603,-15948,-21141,-14909,-14690,-11717,-6598,-15305,
-3136,-7303,-7705,-23711,-6717,-12024,-16381,-21245,-31088,-11533,-11269,-7860,-5897,-9768,-12416,-13056,-4465,-12570,-11543,-10298,
-8848,-10781,-6709,-10051,-10001,-9706,-6222,-20117,-30069,-11123,-21183,-12409,-9212,-7559,-9698,-13912,-697,-6717,-3319,-15756,
-22249,-22407,-3605,-18205,-7351,-7732,-16097,-8661,-25680,-7172,-22241,-15961,-6352,-7570,-16729,-13865,-952,-14071,-5154,-7873,
-28092,-31480,-8496,-16383,-10404,-4734,-22377,-1683,-49468,-7596,-19655,-2062,-876,-11681,-14839,-13160,-3467,-6027,-8708,-4022,
-40599,-45059,-12302,-9975,-5616,-13102,-23924,2899,-48041,-5715,-22493,-4538,-4069,-2895,-13175,-16505,-1867,-3571,-6087,-363,
-45302,-52354,-9452,-1729,-5108,-8921,-34095,-817,-54442,3279,-26970,-1655,-13097,-7432,-7694,-8676,-1405,3298,-5966,-1857,
-44303,-47309,-4282,-4465,-13265,-13499,-13361,-3419,-38944,5411,-36695,-2223,-10611,-523,-19485,-14956,2567,374,-5176,-2919,
-61465,-57468,-9630,-3462,-15401,-5676,-50967,13242,-65050,4445,-33500,-2427,-12020,1953,-17079,-7561,-472,-7016,-11396,3727,
-59211,-45174,-2989,-6727,-16612,-21356,-46312,6148,-56514,13165,-35521,-1591,-7147,-3887,-11325,-5847,-1304,-2812,-8630,-17,
-31637,-38389,-11761,-3276,-27279,-26547,-26777,10210,-26016,3069,-44344,-5175,-6512,1793,-17864,-13285,5884,189,-13683,4342,
-17008,-28877,-8502,-8377,-32526,-18626,-42436,4972,-26551,10785,-48135,-12641,-15313,3209,-13420,-8707,3191,5037,-18878,-224,
-28908,-14703,-9991,-12931,-34968,-23590,-54475,8144,-34159,4745,-45410,-10818,-16959,-1625,-8804,-8453,-5093,-4972,-8197,16982,
-27625,-6021,-1763,-15244,-42674,-30990,-20512,6753,-10067,5597,-55272,-5901,-20191,-3816,-24397,-7303,3787,-9150,-18438,5970,
-20389,-471,-13064,-16880,-38454,-22805,-13983,-2017,-19704,9834,-51025,-19384,-9088,-6046,-18428,-11384,1604,-2123,-28076,8021,
-38633,7061,-10412,-4353,-33474,-19023,-6586,-1583,-15019,8333,-35281,-11925,-19543,2844,-24498,-19897,-7055,-1754,-24574,-3224,
-29424,2102,-12354,-7652,-20566,-24342,-12191,-1491,-20844,3378,-37122,-20124,-17277,2251,-7783,-12200,-10656,-7293,-22315,4238,
-30691,-9615,-9985,-5477,-22669,-23097,-4333,-16482,-5723,-7112,-25338,-20586,-16363,-12909,-17308,-14407,-20658,-6957,-19567,-1345,
-27402,-5554,-20114,-15707,-12311,-21601,-11862,-34083,-9771,-11219,-20565,-33285,-5510,-10103,-14504,-13255,-39756,-15324,-24095,-18283,
-23759,-9332,-12120,-14695,-20794,-16714,-10278,-41276,-12415,-17194,-22794,-30649,-10095,-5671,-15553,-15833,-36583,-8866,-26282,-18552,
-25406,-16084,-17854,-16054,-13758,-23661,-4448,-34427,-6617,-10222,-18907,-21644,-13830,-8887,-20961,-12069,-41136,-8739,-26223,-12489,
-22687,-16441,-9025,-13217,-19662,-24934,105,-38893,-7183,-20000,-17028,-22964,-16912,-9756,-21051,-7200,-34334,-14794,-22071,-17599,
-10017,-12802,-12696,-14588,-16427,-20128,-1033,-13995,-14474,-8725,-11812,-13578,-8236,-8106,-11668,-13296,-35618,-5467,-27711,-12816,
-23071,-2986,-15410,-15100,-13475,-21346,-13626,-18421,-17068,-3019,-16918,-15351,-6590,-10574,-12667,-3534,-29897,-10916,-25534,-2225,
-26350,-2706,-13910,-5073,-18835,-24986,-9610,-14759,-16086,-10432,-238,-23889,-8881,-7373,-15747,-3227,-25405,-3623,-20543,-5269,
-17881,-6987,-10881,-17833,-18890,-11986,-2605,-12384,-13523,-4469,-3660,-26594,-18333,-6976,-17300,-16854,-14833,-7770,-10771,-211,
-9401,-1719,-19840,-19174,-7029,-14131,-9653,-13324,-10036,-322,-3038,-16521,-6033,-12832,-26434,-16033,-7026,-3663,-20639,-13893,
3287,-8498,-14182,-26983,-8473,-9621,-5997,-20493,-27039,-6846,-21178,-15304,-5627,-12952,-5396,-6692,-2593,-11576,-7907,-456,
6702,-11060,-1180,-27468,-11256,-12371,-17826,-15993,-32883,-7832,-22698,-9173,-4793,-8043,3634,-14062,-6767,-12675,909,-7465,
5625,-18176,-910,-20123,-10773,-466,-9188,-8774,-32634,-12027,-33277,-14557,-11875,-9644,-542,-9943,1709,-10385,-413,-11001,
-2031,-22650,-15562,-20151,-2309,-9926,-8855,-3166,-33057,-9622,-30464,-8886,-703,-16280,1129,-7931,1842,-3312,807,-7054,
-4113,-39890,-8461,-24170,-1554,2565,-19206,2813,-36625,-10686,-35985,-10175,-6213,-7137,9401,-11409,4193,-5705,-6751,-7143,
-8750,-41388,-11345,-14783,-8538,-5272,-15190,-1754,-35221,-3691,-40151,-12094,-2666,-5023,11313,-15157,5187,-4215,5425,-8570,
-9918,-51685,-8085,-14664,-4147,-5547,-4446,-3760,-35091,-185,-36260,-3455,-8376,-7323,25685,-5319,6915,-222,-5272,-2974,
-10490,-62236,-8703,-8337,-11369,-708,-16197,12581,-35549,1920,-33022,779,264,-1579,35586,-14587,1607,-7406,-4118,-5548,
204,-66618,-746,-6034,-7669,-6548,-17084,10967,-36011,4328,-40453,-12440,-8490,130,30304,-6458,2940,-6938,-1735,-987,
3906,-59644,-3838,-1198,-22595,-8263,-28772,2713,-32419,10691,-42139,1172,-1428,-4142,29650,-11547,4317,-3393,-4590,-618,
5748,-53462,-8231,-2599,-25723,-13190,-34686,6500,-26852,8845,-41154,-4638,-6683,3398,30399,-7098,4440,2818,-4685,-756,
8900,-42863,274,-4207,-24535,-12500,-45379,12070,-20555,1478,-40966,-1823,-12965,8247,25474,-5726,6013,-7121,-12532,8254,
5386,-29951,-10477,-469,-21934,-17679,-53515,10953,-15722,16852,-39314,1691,-9931,-4275,23490,-14146,-1555,4331,-17049,2713,
10448,-18040,-5758,-9811,-29487,-20229,-46070,12418,-6693,4423,-44566,-4259,-12306,3774,12329,-11269,1861,-5737,-14292,11178,
15144,-11790,-1843,-6282,-35088,-22804,-35169,6197,-10031,14034,-47007,-6549,-19246,252,8239,-5849,2121,-4086,-15166,1052,
-2515,-1916,-8941,-12959,-39917,-20238,-19087,7280,-11117,7987,-42555,-11087,-12215,-7159,-8733,-12091,286,1120,-23685,7579,
-18882,5727,-12878,-2852,-45066,-32635,-17865,3838,-11246,3068,-48611,-8568,-12736,-7976,-19224,-11059,1910,-7332,-17862,13306,
-28446,13747,-7999,-9728,-45967,-25794,-18224,1973,-15355,4092,-54390,-18076,-11167,-6834,-20103,-8973,-5180,-3215,-21205,6813,
-34230,7433,-10655,-7896,-32466,-22757,-6837,-4866,-19011,3344,-27120,-10957,-10357,-7804,-16905,-7725,-15763,-1137,-25338,5085,
-15770,-11037,-10758,-7174,-17567,-28469,-5950,-9177,-15044,-7546,-5880,-16614,-4217,-12883,-18562,-3267,-41795,-5371,-27101,-4304,
-28823,-14601,-21070,-10386,-15221,-16873,-13146,-32366,-8287,-22605,-20167,-20958,-15317,-8448,-22649,-3813,-39019,-10556,-29834,-13408,
-27675,-14493,-12617,-12299,-10960,-13900,-11287,-34813,-16162,-17766,-16710,-29929,-7019,-16104,-13048,-15511,-41231,-13614,-24781,-6251,
-22809,-6322,-15185,-5835,-17477,-27412,-3451,-14964,-4245,-18143,-16929,-14002,-17051,-10200,-22847,-5416,-34829,-15854,-28043,-4408,
-7558,-3220,-13715,-3832,-11668,-24866,-2771,-20521,-11289,-14945,-11210,-12286,-11637,-6747,-8632,-2355,-30318,-16601,-30911,-8958,
-17439,-3635,-13891,-8398,-18411,-21490,-10500,-8039,-12490,-371,-6215,-21181,-10016,-2255,-9777,-2872,-21755,-10090,-29391,-2372,
-5377,-11456,-5613,-5986,-7585,-21821,-1097,-16435,-12317,-7598,5078,-21040,-16115,-7520,-21118,-4963,-13983,-1830,-22347,-12390,
-1441,-5101,-5621,-20125,-8646,-6875,-14096,-10398,-22882,-8405,-8924,-17650,-7583,-17720,-8263,-7173,-10008,-3221,-11684,-7399,
-1828,-5685,-15500,-17664,-2654,-12882,-6388,-8663,-22027,-12307,-18956,-6254,-3657,-11193,-7111,-12896,-194,-6745,-9635,-14473,
-2768,-10694,-11736,-29366,-1305,-3881,-16750,-2098,-27631,-14750,-35249,-12127,-10344,-10535,-2049,-13890,-659,-8531,-111,-18271,
-6141,-18913,-6269,-20800,6463,-4349,-10141,-6810,-32644,-13033,-33795,-9342,-7979,-12860,-869,-5918,2911,-11809,-1855,-13536,
-4965,-31998,3881,-27637,2186,2406,-21500,-9046,-38037,-13381,-26588,-1473,-2763,-11272,13453,-4180,1013,-2631,-5637,-17348,
-13446,-36015,2262,-18076,-3477,-4666,-6408,-4088,-30596,-16894,-33381,-775,-10061,-553,21405,-1661,6783,-8596,5173,-20237,
-36523,-43539,246,-10492,5464,5028,16136,483,-28577,-4368,-24230,-7907,-10130,-4016,34362,-2728,1476,-5071,-5,-20193,
-48781,-48230,-3590,-15915,-1030,-5316,20326,-11202,-26003,-12225,-21211,-6430,-933,6869,39891,-3557,9573,3939,3667,-13699,
-54422,-45242,-5654,-9854,-8011,-3701,20841,-1558,-23853,-9279,-24534,-5071,-1793,2228,42612,-595,13247,1482,3418,-18790,
-55462,-48668,820,-9208,2082,-3358,15019,-3178,-26111,-6910,-21103,3858,-9041,1295,51943,-2130,13656,-891,-8821,-4587,
-45785,-48336,-10445,-523,4616,-9458,3531,-1976,-22876,-616,-26424,-6625,1661,4352,52205,-6971,17480,-4970,-7874,662,
-30396,-44511,-5193,8063,-6817,-7538,-7994,2640,-18533,-1318,-30109,382,-3322,-2318,47725,-5823,18587,-12303,-8472,6458,
-19518,-34872,-1615,6068,-6297,-16855,-22924,2731,-14058,5039,-25403,-4439,-1999,-7060,43381,-2420,16581,-750,-11192,-14,
-9129,-26764,-1459,-3543,-16644,-12870,-32112,2823,-11329,5677,-16883,240,-6601,-1015,40513,-6472,7352,963,-11545,6306,
74,-13629,-6390,-4422,-13898,-17042,-37942,3887,-9674,5342,-20502,3258,-15019,10713,34453,-10730,5628,-4678,-1165,7545,
3820,-3993,-6825,-12881,-14613,-16489,-30901,10653,-5625,12075,-17126,-5280,-6315,4723,23164,-9318,-303,-5939,-8932,3774,
7268,1009,-4171,-5336,-24211,-13294,-30011,2334,-6176,10265,-18230,-10009,-12954,2621,20667,-3415,3089,3665,-16454,-1211,
13216,6140,-7869,-9584,-26104,-16784,-19171,4416,-6654,6596,-18248,-6752,-8339,-1369,9952,-3344,-2485,-2218,-12310,9709,
13546,5419,-8148,-5766,-28894,-21806,-17575,2137,-10901,13069,-19473,-7877,-11852,-1478,1044,-9047,-11572,3979,-10234,6788,
2521,7553,-6118,-5281,-39212,-24063,-7699,3889,-9076,5844,-44619,-12612,-2959,1299,-16670,-15413,1788,1282,-28976,-3354,
-14759,8053,-5171,-4937,-43532,-31967,-11927,8409,-10720,508,-45513,-12720,-12817,1699,-18359,-12025,-8107,-6137,-21428,4496,
-32653,7394,-13870,-929,-30302,-25877,-2097,-1362,-12001,5582,-28726,-13609,-16765,-408,-17985,-10123,-18234,-5726,-21932,-1774,
-22437,-13139,-17746,-5855,-14156,-18819,-11301,-14126,-9452,-9106,-9813,-20386,-5082,-3519,-22508,-3331,-37604,-16152,-31315,-6968,
-18562,-8071,-15409,-6316,-19465,-14551,-471,-21867,-14048,-16957,-13454,-22312,-10343,-2974,-21857,-4716,-38706,-15022,-32581,-12443,
-21352,-14027,-17261,-10644,-10645,-17490,-11124,-23613,-10975,-18281,-15229,-27728,-12882,-4152,-16800,-13182,-39375,-10808,-26599,-7011,
-10827,-7622,-10171,-4584,-20764,-22216,-5159,-22240,-14818,-3646,-27741,-23839,-15607,-7196,-5506,-8912,-23627,-7952,-18397,-7876,
-88,-11275,-5464,-5583,-13009,-19834,-10878,-14058,-8934,-12005,-9812,-21974,-12185,-3858,-12988,-13025,-14792,-3006,-22528,-8775,
-3908,235,-5917,-13016,-11398,-3820,-4545,-13542,-17992,-16515,-17391,-14872,-13907,-14236,-8451,-11410,-13623,-12352,-3401,-9556,
-1150,-13213,-5633,-15545,-143,-2985,-3436,-11468,-22089,-16524,-20448,-12203,-11920,-11391,-9306,-7770,-10683,-11720,-620,-11034,
-3690,-7831,-8659,-30400,2783,-3473,-13453,-15157,-20880,-23422,-27680,-5953,-4811,-13664,-5145,-9259,-2774,-719,-3869,-17939,
-1174,-4942,1604,-28686,-127,4673,-8554,-9020,-27306,-22376,-28759,-11327,-5365,-10968,-565,-2569,-5780,-2097,3099,-23681,
-7511,-10367,-689,-21342,2390,2822,-4836,-1302,-27233,-24442,-26617,-384,2734,-10326,-1407,-5839,-2420,-9555,2584,-16424,
-22170,-9791,2446,-18996,10973,1239,3554,-3338,-28708,-18977,-20213,-9545,4975,217,7976,-3810,-4501,-9403,6981,-18607,
-30071,-13291,-8825,-11459,8006,8578,11405,-4396,-26843,-19217,-21799,-3368,-1787,4099,15319,-3193,2953,-2798,4480,-18994,
-43046,-13897,-3096,-5041,8551,715,15181,-7060,-27288,-19949,-16002,-5207,5664,-4494,25224,-5128,5141,1216,4437,-12438,
-63297,-14835,-330,-8058,10608,9477,14629,-7393,-25901,-11170,-15082,-3589,77,9443,35003,-4752,5521,-7164,5217,-13953,
-60974,-20524,5997,-3012,13109,-1597,15192,-12041,-27563,-11881,-17731,-7785,-4151,6986,41783,2924,12574,-828,5687,-11616,
-50523,-22765,165,-3779,5490,-5539,11334,-7815,-25540,-9922,-14811,4869,4595,337,43862,2173,17312,-650,-3066,-8333,
-37776,-23133,-8163,8030,2751,-284,-1419,3633,-23345,-2750,-20926,4383,2713,3396,42554,3701,21195,-13490,-6832,-10109,
-25094,-19631,-6520,6953,294,-7710,-10781,8270,-18507,-1669,-18387,-517,-2458,-1774,39723,6904,17630,-8346,-3491,-5552,
-11718,-15258,-8706,10318,1477,-11238,-23770,4523,-12460,1450,-13522,-2988,-2170,-3809,30227,4411,15584,-3461,-5787,1523,
2443,-10905,-7372,4296,-11447,-5504,-29916,1385,-8692,4224,-4327,-2394,-424,2731,25914,-4816,5547,-1704,-1866,6712,
11236,-4128,-9657,-6212,-12157,-9668,-28811,6273,-5386,1023,2539,3398,-2724,3401,16542,-7917,1047,4658,-5519,10987,
2616,2958,-11154,-1140,-11515,-8903,-27655,11139,-4460,10320,2497,-5340,-7935,-296,17860,-9692,-7138,6609,-1483,3911,
6978,4353,-6129,-200,-17296,-11867,-21496,8229,-3685,12241,-4709,-3298,-14930,8313,10966,-1752,-3022,-7234,-1336,424,
17376,8690,-921,3849,-27233,-23971,-18586,9811,-3510,2274,-5970,-8223,-3251,-389,1511,-3879,-1378,-6778,-7428,3444,
5969,10363,-9671,5635,-19029,-11694,-14544,4846,-10120,9678,-11956,-7000,-4629,-1638,-9480,-3502,-3635,-4190,-16208,5091,
1036,8627,-2619,6900,-20804,-24386,-15114,8029,-16482,2781,-19324,-7393,-6236,-3042,-23935,-9614,-10808,228,-14763,9142,
-6642,3007,-9254,-3771,-34078,-26148,-6444,13922,-19641,1509,-41733,-7232,-14344,1445,-30558,-5716,-11960,4280,-18901,4402,
-14175,10000,-6297,-3871,-21442,-24386,-6991,-693,-23406,10358,-32255,-8975,-5158,-4915,-15136,-6638,-18361,2470,-29359,3063,
-23046,-11705,-10281,-3425,-15540,-23296,-11800,-13752,-6814,-3295,-16825,-15373,-10070,-6744,-26467,-2461,-35279,-10300,-31890,-11271,
-31935,-16769,-18863,-15529,-23528,-16404,-12650,-43154,-5993,-21544,-17938,-22328,-11523,-15982,-20415,-2674,-32211,-13947,-26552,-17569,
-27156,-10916,-23153,-13040,-20506,-20239,-5140,-11751,-2897,-8176,-13141,-20685,-12159,-12533,-15563,-12075,-34023,-6076,-25740,-4910,
-3899,-2629,-9850,-7860,-16597,-17887,1785,-9230,-9132,-6457,-30929,-12663,-13814,-9969,-8865,-7599,-24654,-7073,-21600,-3000,
-5754,-8997,-9475,-11354,-3862,-17153,-8949,-13142,-5733,-6943,-15576,-22235,-9505,-5679,-17705,-14594,-21566,-10055,-4755,-16005,
-1036,6142,-2714,-15477,-1926,-6191,-46,-12524,-6888,-8399,-3512,-4956,-12454,-13371,-22783,-5721,-16073,-3771,-11630,-6378,
-4961,9393,-4299,-13619,8146,-8731,10292,-17825,-15127,-12235,-9257,-9800,3912,-6181,-18172,-1504,-9935,-12168,-5981,-12406,
3552,21563,479,-4513,4439,4635,25818,-10945,-20292,-29446,-17179,-7083,2262,-12485,-19215,-10159,-9587,-2756,-610,-12816,
-666,22504,2055,-11019,-151,4763,28414,-8309,-18021,-26499,-21050,-7573,1780,-6384,-20940,-4609,-4840,-11290,5827,-18844,
-10953,24080,-744,-13464,11118,6247,31035,-3119,-20399,-26219,-15753,-975,-176,-7996,-18182,-6788,-7078,-7351,6223,-14079,
-18096,18832,-1847,-9879,16625,2695,24298,-12579,-21209,-21348,-9943,2571,6840,-5947,-17595,-7851,-1373,-69,2492,-13837,
-28267,11106,-7530,-4228,11648,14035,20439,-1011,-23500,-21296,-7966,-789,37,-5012,-3227,-2500,-3672,-1646,10872,-10835,
-34717,3710,-8024,-553,21267,1201,14942,-1962,-20680,-12663,-3854,-4915,8212,-2162,2934,-5809,3172,2202,706,-14593,
-46690,-4032,-802,-266,13917,6688,11012,-6163,-18837,-1556,-4795,-2120,-2606,1862,11986,5871,3158,-7044,7110,-13014,
-46011,-10814,-6292,3459,13482,2148,8389,-9751,-16065,150,-5163,-1024,-3029,5896,17714,4523,9945,1179,3309,-12051,
-41980,-13656,-7831,2618,9459,5664,4893,-5475,-13193,-1169,-6040,-6813,3503,7784,20781,7632,14838,-8439,-2352,-3153,
-27766,-11192,-6474,2044,4965,-499,-416,-219,-10268,-3792,-245,3357,2169,1799,22231,2819,13240,-2892,-6974,979,
-12075,-4566,-3677,6597,-4729,-1013,-5806,12203,-6490,948,153,-719,5206,-9915,17165,3652,6061,-6764,4349,-2076,
7662,-2015,2836,8401,-5134,-3552,-12310,6011,-4196,974,-335,6623,-9946,-6322,8644,4699,6080,-6370,3814,2501,
18542,-3686,-4391,-3410,-2360,-6531,-15044,6492,-2230,5242,10371,5583,-5555,4978,2770,-4033,-507,-799,-2283,6465,
25902,-841,4115,-4305,-8891,-10699,-17435,4909,-1703,2746,12476,-2782,-6994,1189,-899,-1725,-200,8171,-5657,4099,
18672,2620,947,-4470,-10406,-16029,-19647,10891,-296,1964,11303,2923,-9566,6762,-923,-1706,-588,-3040,-2735,7032,
13273,11031,-2436,-3645,-13806,-13077,-21480,5927,681,11952,7921,-6501,-8581,3462,-3819,1948,-836,-2598,-10579,-386,
18974,8014,-9741,182,-15184,-22550,-16558,12773,-3619,11794,9588,5996,-3573,-3570,-9818,-5283,-8904,-3088,-5059,7673,
18950,7400,-143,1319,-24824,-13853,-16989,3817,-9833,10869,7773,-1567,-7944,1912,-28124,-4233,-10085,1286,-14146,2738,
6439,7561,-7894,-3245,-23743,-20567,-10840,4615,-18233,3376,-14876,2278,-1059,6053,-41378,917,-5613,-7424,-16059,7113,
1442,2700,-3752,-2598,-25784,-29709,-13075,7964,-21469,7646,-26148,-5149,-6641,2299,-26316,1278,-15734,-4532,-17835,7542,
-11624,14522,-3629,-1615,-25108,-24919,-5592,1886,-21913,4380,-39332,-13420,-10576,-4715,-23145,-3094,-16863,-1449,-20652,5178,
-31640,622,-1046,-6864,-29827,-18720,-6001,701,-6279,894,-17028,-14755,-6095,-1965,-24831,-4477,-24811,-8333,-31065,26,
-24953,-13593,-13567,-4294,-11657,-9825,-11241,-53999,-14817,-28827,-22503,-41847,-17770,-10504,-9319,-12394,-31624,-19243,-25008,-20202,
-27209,717,-10918,-10412,-15940,-16365,1976,-17988,-6785,-5588,-24227,-13058,-5740,-8682,-19965,-9918,-27130,-8797,-26143,-320,
-25420,-4489,-7773,-3512,-10183,-8345,5457,-22932,-3655,-13399,-33908,-13386,-5633,710,-20547,-5295,-40830,-13269,-16673,-6081,
-4697,8015,-11746,-2997,-3857,-7459,15384,-17266,-7241,-6696,-6414,-12856,3143,-10855,-27219,-10219,-35252,-166,-8055,-6118,
2849,19998,-12194,-2740,-1909,3604,19317,-11000,-4243,-19411,340,-4406,-3968,-6912,-38271,-8442,-17926,-5812,-12375,-7270,
3383,28462,-3258,-7219,4910,5026,28953,-16452,-5414,-13851,-145,-2783,-5673,-12993,-41837,-8081,-17132,-2027,-5670,-15852,
3219,33412,-8692,-5264,13200,-765,30222,-16376,-14280,-23668,-4430,-10672,948,-11102,-37896,406,-13671,-208,1341,-13386,
1009,28519,714,-5068,17289,4626,36318,-12440,-12897,-23418,-8305,-4512,-3866,-6154,-39184,-7727,-10686,-9191,3560,-11914,
-2986,29459,-30,-6915,9194,9633,31327,-14343,-11507,-19514,-601,-5390,2101,-10056,-34028,-9051,-11096,-502,7696,-13918,
-8900,20541,-5481,-4873,21075,5988,26575,-6410,-11144,-19101,240,-2096,-766,-7608,-35692,-3936,-1654,2033,1127,-12514,
-25877,13848,-7395,-631,19826,1657,14873,-7664,-7476,-4328,6991,-9007,3956,-1422,-29096,-6231,-3588,2704,6956,-14849,
-27914,458,-1846,-1919,12988,4411,10345,2423,-6394,-8232,14751,-1597,2373,-7071,-16985,-1598,-3859,808,-951,-1129,
-30902,-8679,-6965,1,8830,-2190,3723,-6679,-3257,1944,13336,-6485,4807,4573,-10409,4499,1501,-2160,2333,-108,
-32588,-11355,-6082,6105,4059,-3520,324,-4252,938,5474,15624,5033,971,4430,375,-5021,2651,4977,-279,-4068,
-34817,-8164,-4611,2704,-1240,-3630,-1635,-2719,4984,1557,10421,-3210,-794,6125,5940,2810,5903,-7171,3128,6537,
-20448,-1286,3784,377,3382,-5218,-3177,-2462,6656,1056,8981,-3111,-1516,2271,3285,2241,7403,-8978,-4384,7561,
5576,4451,-4827,5477,-3709,-10830,-4756,3918,6662,-1092,6083,5555,1792,-3471,-5383,-783,6309,-4290,4634,1441,
26428,4967,-2789,1377,-2765,-8066,-5599,14388,4899,-4032,10103,-4205,-5027,-1434,-10799,347,631,2015,3366,-1814,
33557,1070,2065,-6287,-1031,-2720,-4505,11451,2025,-1233,17308,-513,-4009,5074,-15207,-2153,-2667,-3586,-2422,6137,
35071,288,-422,-1553,-9653,-8553,-3360,8581,946,-242,14882,850,-10263,6275,-15341,-3130,-861,-328,2867,5269,
25643,5866,-7994,-1633,-10399,-13014,-8429,1208,2465,10575,17997,6131,-3345,-496,-16592,-651,964,-3004,-4345,8491,
18380,13233,-7941,679,-16430,-14458,-13280,1092,3162,12922,15684,-7942,-5153,5917,-14044,-2450,151,-1844,-3282,638,
25750,12289,-2974,-1270,-23677,-19001,-9509,14911,-3368,5518,17883,-244,-2329,-520,-14705,-6095,-4937,-4130,-5009,2487,
17729,9721,-3181,7889,-19343,-14767,-13375,2215,-9131,2181,14889,-3509,-13374,48,-38078,-9145,-6323,5692,-14794,12620,
21976,2258,-295,-3714,-26932,-21980,-10784,10127,-21231,2405,8152,-8339,-2778,3041,-30407,581,-10603,2986,-22055,5427,
493,5266,-10141,7168,-25956,-26016,-15428,10100,-22241,8594,-27117,5115,-13663,481,-32033,2476,-12587,-2228,-20088,1796,
-8152,13393,-2660,-1712,-27850,-17151,-8687,3864,-19749,6561,-34337,-2855,-13057,794,-21443,-13490,-20288,2874,-28953,348,
-30979,5682,-1430,-3547,-21131,-27448,3912,-12006,-16602,-1996,-35923,-15030,-12748,3694,-18169,-12188,-22285,-2858,-22713,5035,
-30619,-16380,-20065,-2796,-13773,-15062,-5380,-25943,-2744,-16489,-12787,-22153,-11887,-16588,-23901,-9740,-36791,-9242,-26718,-17474,
-21080,-9685,-8824,-4968,-13875,-13555,-6205,-24776,2180,-12583,-27460,-10598,-13175,-5734,-23700,-12248,-39198,-5711,-19966,-4012,
-26313,-526,-8811,-3710,-7254,-11341,-3241,-14621,2898,-3372,-31006,-4388,-3551,-9367,-34504,2705,-50277,-11989,-17255,-2283,
4677,13374,-11355,-221,-3042,-6343,11801,-16961,1196,-12247,-2666,-11171,-6307,3102,-49262,-2907,-35582,-8222,-6119,-10634,
6930,11064,-15265,1239,9475,-1499,21935,-15418,-5081,-10631,10729,-13628,-3462,-5940,-47547,-3075,-31692,-3867,-2993,-5627,
8238,24241,-2585,3267,9603,7773,28185,-20636,-6441,-15730,9912,-1718,-3213,-7644,-51296,-6850,-24662,-10100,-4498,-12775,
19887,25264,888,-567,13815,2905,34304,-22878,-10923,-25527,5228,-8433,90,-5741,-50102,-4972,-17224,-2906,-1141,-12183,
8790,31891,-2081,-8747,10054,736,31684,-24134,-593,-19752,7261,-4678,-1463,-6303,-53652,-6392,-11982,-8175,5800,-5714,
7338,27694,-1654,-7386,7608,6600,28469,-13069,-1021,-17732,14073,-1566,-612,-6098,-49988,-7009,-9298,-2402,5667,-14374,
-14205,19054,-2903,1076,12623,7816,17847,-10506,3246,-6860,14426,-7126,-277,-6495,-52772,-3467,-2391,-4794,1833,-11313,
-23119,5179,-8176,4504,7635,-1735,10372,3129,3256,-6201,15920,-7140,153,-53,-47501,3102,572,-5705,6855,-10928,
-18827,-11442,415,3515,2640,-635,8857,3872,3885,-1303,21215,3628,-5223,-1626,-36819,2530,-482,-3833,-4035,289,
-15421,-16660,-2115,-1348,-9642,-5517,4999,-804,8814,1416,22498,-2117,-1360,2542,-21514,3413,-1905,2356,6217,8610,
-17004,-11344,7194,-3221,-14103,-10500,4017,-861,12322,4381,20035,-3558,-3870,-733,-8734,2629,812,7975,2739,1097,
-30572,1628,859,-2145,-7351,-10494,936,-6378,17739,4816,12873,-6153,-8749,631,-6,-2804,1853,4850,4211,7924,
-17348,11815,-186,-3440,487,-12155,-361,5462,17787,-1289,8549,-3027,-2758,-5004,-4812,-630,3992,-5409,-132,7509,
8596,16358,-10487,-2627,-1840,-3447,-2663,12175,18084,76,4896,-6253,-1523,-13039,-20234,4623,1326,-4104,-181,4883,
33672,9757,-4720,-11236,7518,-10765,-859,13690,13926,2568,12777,1601,536,-5896,-30956,898,-3040,1453,-5378,-712,
35453,2877,-4042,-9033,2285,250,3040,9009,6018,3627,18403,3342,-2634,-1055,-28167,-4195,-8547,1385,-3582,6536,
43426,3711,5392,-1491,-7025,-1306,4121,5577,1529,-612,16390,-5034,-3933,-32,-28540,-903,1204,397,-8033,1852,
31719,10883,-6937,5909,-17557,-11950,-1578,6186,3800,3062,19155,-6169,-8226,-1875,-25115,-1822,-553,-2929,5439,5428,
28572,15815,-3827,100,-19673,-16878,-5369,9070,4368,6549,26835,-2110,-8054,1692,-28084,-7162,-955,-564,-3491,-663,
26756,16783,-9893,9475,-24988,-11825,-6298,11111,-935,10556,22698,1252,-15123,-6210,-31172,-7496,-3064,2328,-5514,-2759,
14571,13519,-4070,7333,-22563,-28787,-8743,9300,-10064,2513,21828,-11040,-3778,2527,-30644,-5914,758,-2188,-15763,-794,
-1822,10545,-6936,4923,-20246,-23844,-10771,6415,-21749,6730,17016,-5995,-3817,2067,-34438,-796,-7945,-8880,-18228,7535,
-10749,14252,-13596,-1821,-16819,-13592,-14046,4835,-24188,8634,-29642,-3189,-6928,7297,-31079,-10465,-20461,1309,-20510,8305,
-17092,11780,-10358,-4933,-37086,-26498,-543,4807,-16727,4844,-52590,-5016,-9703,67,-31619,-8109,-14324,2435,-20212,717,
-29284,7738,-15984,1757,-26497,-17636,-4260,-9477,-6462,338,-25682,-13414,-13018,-1239,-24526,-7738,-24996,-3101,-26163,-1412,
-27821,-6188,-19197,-13343,-22658,-16300,-5883,-20398,-3510,-15440,-13145,-17692,-13417,-4132,-23412,-5210,-42713,-4359,-23682,-11826,
-11692,-10237,-11239,165,-3896,-20090,1060,-10530,-7827,-9383,-29818,-6635,-10793,-5970,-17257,400,-48021,-9832,-12397,-8155,
-20129,-2258,-3964,-974,-6022,-6185,8208,-11626,-3841,-11231,-38088,-4674,-7165,-6612,-38880,3673,-59664,-13160,-10007,-7371,
5922,9777,-2879,11155,-2225,-4540,11755,-19473,-120,-8882,-5664,-9978,-181,-6674,-53562,-7772,-42289,-13160,-11924,-8260,
16665,18081,-3996,-3510,3380,-124,19917,-18004,1904,-14868,17613,-9690,-37,-3915,-59298,-6297,-33506,-8771,-9469,-7740,
25214,22192,-4577,-1242,7096,2898,29084,-19386,-1510,-22013,19572,-7352,512,-4449,-61063,-8457,-28161,-6000,-3546,-9291,
27962,31861,-10110,3,-701,7428,31074,-19775,2941,-19025,17466,-1943,5235,-9257,-67526,-8882,-17594,-13062,2321,-12256,
33178,29533,-9081,2527,4467,6327,29431,-18278,3198,-18360,17109,-15028,-7119,-8234,-68934,-595,-11282,-4953,7257,-13136,
3588,24846,-1784,-1926,8551,2046,20335,-17796,9581,-13474,24977,-5727,-765,-820,-67955,-5543,-2984,-12847,1695,-5449,
-28443,14477,-5788,-987,10390,3565,12626,-3222,10608,-3472,30768,2479,-9891,-5714,-64541,-1372,-4653,-331,-658,-9974,
-41208,-3835,-8782,3606,5997,-6592,11565,-10,8791,2536,27462,-7827,-6227,-5837,-59273,3868,-4154,4853,6417,-3103,
-20494,-19638,-2436,7903,-1830,-2864,11400,13475,7923,260,25381,1565,-9325,-3583,-39332,-4455,-3430,2335,-4201,5565,
-11823,-17135,3592,-2582,-14619,-5696,5578,5042,10015,10265,23151,-438,-4287,-3075,-19043,4940,-3784,-757,-443,8084,
-27553,-4200,49,3753,-11764,-13412,-1127,-133,13634,4041,11462,-8203,-2613,162,-3665,1429,4534,-2550,288,10753,
-31644,10375,394,-4024,-7260,-15963,-2415,-2445,18699,2168,8598,2589,-7242,7742,7372,-9895,5739,3303,-1852,-877,
-22620,20013,-3128,-8249,2958,-6936,-3897,-1355,20777,149,4500,-3665,-6097,-1557,-372,-5024,3683,-712,-4783,6065,
14765,15864,3268,-5443,-676,-14670,-4836,7248,18471,3709,4367,-828,-1484,-12009,-18059,-1946,-4685,-3968,1533,-517,
30062,5047,-4491,-11350,6017,-4694,-1944,5597,12972,3869,5899,2564,-10365,43,-29185,2343,-9462,3232,3224,2829,
37438,-23,-1342,-6906,5968,-4071,3127,4665,5149,2327,9595,-1420,-8860,-1938,-33560,3568,-7784,6566,-2339,4119,
38340,5354,-7875,-2388,366,-5703,7693,10890,2830,7004,12473,206,1267,4092,-36080,-4539,-2052,-3666,-4404,-5112,
36200,12666,-8948,423,-7754,-6839,6042,7863,3080,8435,19090,-10405,-6497,1915,-40681,-1170,484,-2722,-1620,-4062,
32888,19507,-2369,2306,-22452,-7231,1506,4435,7107,2029,27490,-8402,-13950,-1486,-46386,-7331,1186,-1668,-1038,3021,
26856,16862,-1756,2233,-24190,-19171,493,10010,1906,6445,34038,816,-20481,-3081,-25902,-10790,-4481,2090,-2199,-1245,
18423,11998,-1825,6805,-19410,-16957,2348,7809,-10777,10316,27707,-8818,-16455,-2785,-20849,-6525,-1161,-1025,-18307,-3257,
-7838,12060,-12175,9102,-22532,-20321,-6022,4268,-20780,8257,25004,711,-17326,-1162,-31693,-3939,-7994,-465,-15441,5024,
-426,14580,-10914,1719,-27026,-17789,-11119,6150,-24133,4171,-24181,-9677,-2816,800,-23591,-6777,-16171,2148,-19926,5608,
-4301,6069,-7569,-3753,-31982,-24430,1993,-652,-20046,3237,-44772,-14016,-5167,4112,-26570,-4678,-9696,1420,-29634,3967,
-27551,9223,-7693,4089,-31702,-19365,349,-4916,-18577,1456,-32553,-21962,-4990,-2237,-15529,-3120,-23948,-11658,-26652,-2841,
-23301,-1068,-17955,-8425,-18944,-13799,-4898,-19309,-2809,-8875,-15878,-20898,-13221,-8856,-20566,-8043,-38113,-10237,-22094,-3942,
-10262,-6900,-14018,1472,-13812,-11100,-736,-18281,-5364,-17491,-30008,-10479,-3367,-11594,-20143,690,-49815,-6409,-13555,-9497,
-13621,201,-6964,2084,1725,-12382,-5576,-8693,2038,-3435,-41535,-2960,-8494,295,-42191,-2136,-54143,-4232,-19395,-12925,
19029,11290,-4947,3872,-8604,-13154,7353,-17327,1657,-16137,-1126,-5921,-2052,-2051,-54438,-3670,-42835,-4175,-5006,-8118,
31207,18808,-14201,6251,-1668,-515,17817,-17558,7131,-11748,15382,-13335,-7072,-4649,-68565,-8165,-33094,-4809,-3932,-8686,
37930,26101,-4767,-460,-2732,212,23610,-18999,7469,-11691,27342,-7379,-2503,-9086,-76472,-3041,-25164,-16966,-5566,-10408,
35725,28715,-11236,8265,10262,8097,28550,-21038,6706,-8714,27076,-11125,-6042,-11389,-80975,-7142,-18430,-16162,-2147,-7659,
39778,24554,-7279,2821,5739,7149,22957,-19205,8719,-10593,37501,-5346,1094,-10283,-82069,-7151,-7315,-5528,-8763,-10669,
-3597,17957,696,1778,10913,-1513,14648,-9651,12266,-9022,37230,-4069,-7631,-4904,-81592,-2564,-4058,-10699,-212,-3154,
-37533,4593,3111,5943,13198,-4630,12508,5812,11461,1928,33523,-8514,-7665,-9444,-81055,-2933,-3843,-4522,-5009,-9677,
-48588,-11641,3261,395,3760,-4012,12825,6900,6625,7493,27789,-4221,-6512,-3048,-61354,3545,-2184,-2370,-4577,-5188,
-26212,-18849,-3645,8843,-2749,-8476,6868,8631,3698,11503,20042,-362,-7717,-6715,-26622,-2736,-6073,5063,1052,5460,
-21952,-8982,-6057,-1266,-10547,-13403,-3477,4995,5371,6185,12315,7954,-9400,-2656,-3451,5909,-196,5270,-630,9998,
-32343,5023,-1891,2104,-17472,-11324,-8577,-4003,7468,3866,4478,4292,-6397,-107,13725,253,6337,7953,-4761,-2022,
-38038,16555,6317,-5093,-5699,-4795,-4702,-1641,12058,-4240,-2379,-3324,-6414,23,20112,-5527,8155,-2132,-11182,1372,
-16677,16206,-6659,-6175,6361,-6670,-2362,4983,9587,440,-7488,-5321,3148,-8524,7452,2497,5018,-7189,-7916,566,
13069,7949,1147,-13520,4792,69,-4885,8860,9912,-3162,-688,-1404,814,-6785,-9710,-37,-6583,705,-7826,3960,
30503,-1266,6991,-4954,5991,-7303,-3846,7957,7319,2248,79,-4520,4360,-5728,-25794,-1216,-12579,2054,2904,863,
38996,-2482,3483,-1288,3682,-2647,3294,4684,2913,6967,656,3688,-2263,-1815,-36804,1152,-7983,-1213,-1322,-1784,
33446,6745,-7051,-5383,-4636,-1654,9794,-2041,3727,5420,7099,4409,644,1716,-41703,-3898,-3319,-5262,-993,6272,
41926,12490,2563,3400,-10203,-4681,12365,-912,5652,645,12876,1827,-2748,529,-59512,-13467,5685,-8825,-4312,2892,
43254,16736,-7756,6599,-15275,-20031,6015,1983,8031,3719,26951,-143,-13825,-3943,-53881,-6892,7723,-3199,-1658,-357,
28619,14953,-12299,4081,-18828,-16193,6789,11043,4459,2505,34549,-11554,-13361,2875,-31310,-9992,5527,-9196,-9344,1867,
20230,15511,-6269,8331,-22207,-18012,5805,12995,-6923,5260,31888,-14055,-19112,-6419,-15156,-4488,1319,-4974,-13341,-2962,
-5836,18890,-8908,3369,-23776,-26675,76,9328,-16252,695,28819,-10949,-9494,3384,-28243,-6882,493,-4710,-16348,-5269,
-816,8089,-6361,3402,-21803,-19246,-5816,5908,-20418,13392,-10800,-12673,-14365,5899,-19155,-10242,-16958,-3641,-19039,987,
-8429,2480,-3403,-1386,-28123,-25316,-1788,6103,-16902,3634,-37785,-19021,-7442,-4159,-17436,-1833,-16383,-6054,-26943,8070,
-15666,-973,-12540,-8935,-23703,-18309,-3985,-17592,-16409,138,-20980,-11429,-6327,-7822,-7512,-162,-26440,-1659,-22729,-3177,
-19317,-13563,-10681,-7364,-15002,-19016,656,-14330,-10067,-11654,-13904,-22212,-7535,-8389,-18671,-3550,-40254,-16653,-25287,-14870,
-20373,-5072,-10340,520,-4298,-16892,-10435,-22517,-3101,-16154,-34800,-17316,-4397,-3282,-15777,-7520,-43318,-5484,-18088,-8881,
-15128,6132,-7741,2154,-8200,-6192,3696,-19659,-3485,-11756,-47644,-10448,-6251,-1427,-36753,-3788,-53508,589,-11738,-8899,
8598,15244,-1764,-729,-4547,-4496,12171,-20295,5074,-7279,271,-12403,771,-7293,-51020,-8366,-41293,-13903,-14423,389,
38115,16796,-9144,11584,-1825,2287,21442,-16363,2973,-13365,18477,-8219,-7753,-7953,-67259,-5766,-29194,-17247,-9637,-5150,
53272,20885,-6426,1235,-2043,3884,28497,-16553,6152,-8165,24983,-11940,-10624,-9738,-82035,2515,-18792,-17616,-6791,-12482,
51714,25691,-15323,6269,-2210,-1552,19587,-24724,13947,-6821,31300,-11593,-7540,-14948,-93588,1386,-10018,-13119,5144,1426,
36794,22141,-11305,3805,5153,-77,13857,-5093,16043,-5632,42221,-7135,-8337,-10837,-93809,-3658,-8917,-9085,2153,-5007,
-10954,14160,574,5443,9450,-7682,7358,-3640,15477,-5320,43233,-14107,-7325,-5897,-92670,-7971,-5629,-1179,484,-3575,
-50546,-2534,3817,-386,2712,2507,12071,814,10299,2225,33794,-1686,-8268,-3850,-86522,-5242,-5785,-3737,316,1764,
-44745,-13036,5275,1712,368,-12726,9226,10577,3611,7891,22381,3024,-7920,-3184,-46103,-6980,-7217,2680,2614,-2506,
-21210,-14096,709,-1207,-12435,-3835,386,8307,-3564,-13,11483,531,-2326,-1225,-6968,356,-3957,4844,158,10382,
-36214,-1540,-7562,7368,-6401,-4406,-11214,5206,-2835,3230,498,3796,-1407,3871,16056,-6413,-1897,-2820,1743,9877,
-41277,9782,1838,5350,1742,-15377,-9898,-10019,-1490,4619,-8263,1657,3738,-1305,26250,-7202,4983,-3048,-2402,3370,
-38116,16002,4141,1549,1442,-2593,-4009,-9900,18,2266,-17327,-5307,-4469,-2626,34533,-5125,6490,2970,-3779,-9656,
-13686,9094,365,-7130,8398,-2299,-3499,-3597,-1337,-4605,-15346,4153,-969,-4412,21130,121,1562,-2601,-7878,3939,
13401,289,5276,-4760,17755,-4869,-3708,11345,703,-5453,-13775,-5883,-1374,-6795,-4931,1287,-6069,4988,-6804,1085,
24355,-3235,6293,-7650,11622,3645,-2203,9349,2309,-4276,-6964,-325,-796,3623,-22956,-4654,-10332,3126,-9928,3706,
33027,2946,1428,-1203,4370,-8335,5872,13146,4010,-2301,-4455,3747,-183,-4550,-37070,-8047,-10464,2413,1825,1869,
34651,10812,468,-6341,1383,-6934,14609,4795,6730,6499,-574,594,1772,-4789,-58266,-8415,-2353,-8707,-4964,1449,
30296,14626,-173,-9062,-2048,-8245,18067,-3572,11056,7723,10107,-8528,-1662,-115,-64625,-18124,325,-7795,-1014,5802,
36695,17529,-8161,-1234,-9820,-11423,13787,4199,12229,4466,26023,-6763,-12227,-5932,-54609,-14317,6166,-6667,-4511,3884,
32772,17964,-9328,7682,-13384,-14180,8606,1260,8689,4398,36134,-15506,-22463,-3216,-40109,-8523,9598,-2396,-10561,-974,
14507,21758,-12097,7885,-20500,-22787,13374,4502,-879,4518,28046,-11802,-18940,315,-17119,-11491,8190,-15989,-5503,-5337,
-1401,15518,-15088,8232,-23870,-20349,14832,-2852,-18515,-73,23616,-15469,-19806,-7001,-7544,-5458,1928,-102,-4776,2197,
804,7740,-8249,1182,-23124,-27948,-1056,-1740,-14799,10432,1580,-11511,-13303,-6705,-15949,-453,-10607,-2722,-15579,3209,
-9676,10550,-12437,6029,-21332,-15076,5309,-6569,-17316,4330,-37990,-13971,-14275,-5187,-17025,-4608,-10674,-9295,-29051,5893,
-25931,-3268,-18140,-1372,-17591,-20826,-1603,-13971,-1029,-7684,-11756,-20516,-16285,-6378,-15275,-11709,-34023,-9619,-18330,-5456,
-21740,-15827,-13707,-2551,-6513,-23124,-3832,-24298,-10898,-9082,-18157,-25857,-16113,-9725,-13238,-12896,-42541,-10752,-19219,-6099,
-20688,-14120,-17068,-444,-7062,-14129,-8811,-32630,-5161,-19688,-29196,-20255,-8907,-2799,-18471,-733,-35972,-5039,-18176,-8740,
-11213,-628,-5853,-1650,-2073,-16323,2238,-16403,-829,-3763,-27414,-13856,-1220,-849,-35717,-6375,-47126,-11339,-14273,-2950,
19202,11518,-18717,623,-7484,-1519,11955,-15491,-1753,-6163,4135,-9581,-495,-1602,-38648,-4814,-37649,-8548,-11310,-4527,
45039,14594,-6902,-1894,-2745,-11121,19366,-24669,6832,-1569,19479,-7374,-11668,-2709,-68103,-11,-21657,-15502,-7426,-4028,
56262,23531,-7117,921,-1495,-6916,16593,-20568,16683,-5297,25621,-21389,-15024,-10407,-87585,-258,-9024,-10333,-4348,-893,
62244,21541,-13831,6741,-1609,-2259,9435,-11388,16644,-4376,39452,-13060,-9428,-8504,-94034,-5505,-6504,-8678,-5325,-2420,
37766,19854,-5012,2249,2127,-277,4585,-5308,20043,1690,45577,-14174,-12379,-3683,-102065,-4620,-5776,-4532,-2095,-9161,
-21864,10255,-6255,-3223,6659,-1784,6194,450,18532,34,39881,-9228,-6023,-5278,-103320,-6914,-4406,-4371,-2171,4076,
-42141,-3646,-5926,-1407,-2256,-2189,8247,-5051,10794,6690,23718,-6463,1397,-3815,-87857,-6893,-1440,4855,1087,1560,
-24073,-11227,7396,-2541,-5899,-10746,5069,11269,-55,3787,8967,771,3458,-3335,-34943,-2782,-2513,-3967,1219,522,
-15651,-7066,3649,-2252,-5677,-4106,-6446,8199,-9395,1543,-795,1984,-2254,-1721,1453,2829,-3439,2180,-3443,5868,
-28953,3635,-2945,3644,5824,-12049,-16694,7645,-11177,-3525,-8983,8812,6711,6270,22450,-4310,2408,-6062,-4810,3815,
-39245,14093,4414,-4040,3835,-7792,-13729,-1999,-10019,5,-16068,5527,1039,3269,37015,1478,1515,-3993,-599,-6752,
-39514,11869,-6875,-2531,13815,-3431,-4926,810,-9947,-3207,-23805,-3004,5577,-54,43959,-546,2265,-800,-747,-5226,
-9154,5288,5687,3518,15686,-5274,-5692,-4466,-8409,-2801,-24062,-933,605,-2513,26151,-4256,-2419,1273,-1813,-1255,
8699,-2326,-3395,-4037,14726,-513,-780,5968,-5979,106,-18943,773,-2114,956,-273,-55,-10042,5644,235,-256,
27050,-2197,-1690,-2069,2637,787,5040,9339,-2686,-6279,-16729,6940,5903,-3087,-24122,-2973,-8627,-1352,833,7389,
27999,5790,2390,-6897,3840,4388,17218,8086,4357,-1147,-17468,-3591,-1934,-4179,-45591,-6095,-6062,-4802,580,5916,
33564,12688,4177,-9952,356,-7591,20850,8300,11433,510,-9426,1010,-2354,-8102,-65636,-17794,-2305,-5357,1728,3260,
38326,14388,-5472,-14652,1296,-8937,24032,10548,14848,3034,2100,-2023,-10460,-7187,-68802,-21827,3489,2273,-5556,-1304,
25056,15935,-11863,-10701,-11384,-8673,20520,5252,16449,1198,24019,-10277,-9632,-2978,-52608,-24583,3536,-6668,610,8269,
31998,20752,-8661,1416,-27612,-14372,11165,-1037,11589,-834,40288,-14406,-14961,-9336,-46578,-11199,7074,-5345,-336,2104,
19963,19190,-11182,15525,-19588,-15240,18069,-7200,-1613,638,22530,-21066,-25289,-5985,-23452,-7013,14409,-13714,-6353,-2135,
6284,15798,-10054,7808,-27220,-18248,10456,-5227,-7930,-12604,17110,-21767,-13028,-1635,-21429,-2532,15991,-10327,-13275,-825,
-2851,4468,-9890,4348,-24850,-25114,415,-7609,-13939,-5518,11271,-5931,-5575,3320,-18087,-13821,-2171,274,-19700,169,
-43181,6658,-13943,-6185,-21342,-25619,1813,1138,-9415,-1044,-30957,-16431,-8406,2230,-20875,-11322,-14546,-5164,-18361,366,
-15180,-7353,-4497,-10054,-26183,-25804,-850,-10344,-2197,-12295,-10923,-10138,-7355,-3053,-22324,-7195,-33930,-6410,-29968,-1593,
-10713,-5541,-19302,-10338,-18468,-21576,319,-16916,-12592,-12041,-17143,-11942,-16403,-5370,-12801,-1466,-42663,-8998,-31994,-6664,
-9882,-2562,-10590,1618,-13291,-13101,-8987,-37248,-10500,-19064,-27719,-25157,-6577,-9901,-13688,-11274,-29894,-6922,-22915,-15083,
-2349,-1664,-14910,-9319,-7967,-12329,3400,-16360,1547,-10254,-21605,-10209,-4922,101,-36980,-2313,-32586,-11789,-21138,-5421,
27036,4874,-14299,-75,-10617,-2950,13931,-25091,-5950,-10259,220,-7057,-4241,-1343,-35551,-5763,-30169,-7369,-15026,2521,
38127,15357,-8159,1480,-7886,-1614,23670,-15124,12174,-7305,15110,-23745,-16116,-9950,-59101,-10857,-15816,-13490,-4261,5442,
46509,18832,-16624,3841,-5877,1636,13235,-16172,21925,4851,22479,-19308,-19303,-7205,-84039,-4931,-4234,-18301,-3021,5251,
61252,17654,-13525,9680,-6819,-1705,1527,-6645,20504,421,37272,-12139,-14342,-7198,-97598,-2256,-3589,-17653,-1450,6236,
37969,17024,-4662,141,-3815,-4744,-202,2817,22232,5567,44371,-15202,-13583,-8329,-104493,-1439,-6754,-4761,2059,-6844,
-7969,4790,229,-741,-2619,-4098,5935,2639,19153,8980,29288,-9411,-5744,-8537,-107819,-7258,-4235,-8591,2445,-825,
-16633,-5705,1172,-3484,-1836,-3096,6787,3035,10124,7417,12984,-6131,1587,-12974,-83823,-5226,-2406,1325,-3179,5326,
-11024,-7544,1512,3858,-5532,-6788,-2191,12083,119,-783,-3870,727,-2520,-6761,-33134,-5149,-5070,-3324,7418,10573,
-3301,-1983,-1767,-556,-8242,-3356,-12668,5239,-10019,4782,-10888,7808,7858,1094,-3400,1783,-2952,-2884,833,-665,
-16905,9195,5862,10027,-778,-2644,-19826,1760,-13978,-1581,-21454,6553,-2466,-3668,20646,5663,-2801,-4912,4641,-233,
-22006,11158,-5269,1583,6320,-5747,-12373,-10521,-14217,-339,-27111,6468,7110,5697,29917,3145,1866,-4337,458,-2228,
-24480,8171,1973,-3512,14026,-6028,-6843,-5226,-16649,314,-23194,11879,10401,3264,47151,-2605,-4129,1002,-252,-7106,
-7115,1822,357,-4252,12926,3235,-2519,1668,-15699,-3094,-23258,10208,2623,-3285,26250,3187,-6543,6070,-5403,-1307,
12720,-2629,4658,-1661,13196,4274,3368,9199,-8882,-4048,-25849,234,5636,4353,-3964,-4801,-5907,292,-6724,-2334,
24591,-159,-1745,-9515,9066,2632,14350,8951,-2447,-728,-22371,9926,915,-4042,-30803,-3769,-7315,8325,-3012,-587,
20637,5046,-5516,-18679,5869,243,24553,3174,7840,-270,-23022,3299,-1957,989,-58145,-15678,-4695,3218,2302,6014,
22158,10418,-5569,-14857,-1774,-1727,23720,-955,15059,6927,-19209,-3189,-259,-6420,-71411,-19341,386,-5518,6092,5998,
24735,8877,3604,-17318,-3909,-1383,27971,-3115,17587,7504,-4892,-8149,-11439,-1049,-66406,-28836,2570,-5549,2414,3771,
28180,10385,-4432,-8258,-17712,-7125,29232,6429,15457,2157,16650,-5262,-12992,-12383,-51025,-29776,4234,-1822,3296,-839,
24495,11183,-10175,6565,-18396,-18952,19979,-4958,8448,-4196,26801,-22389,-14014,-2656,-48401,-11229,16206,-13074,357,754,
19574,11835,-17551,22886,-12113,-8131,19878,-3991,-319,141,21051,-21422,-25560,-7627,-32831,-11758,13605,-6744,-5058,-7091,
11650,5281,-9199,13451,-24443,-21637,19057,-9596,-6719,-10095,10041,-24070,-11752,922,-32529,-4793,16865,-8034,-2919,-11926,
-3951,-93,-14734,6297,-16702,-20490,8286,-2887,-13856,4421,7456,-17331,-3875,-2035,-18165,-11650,-7421,-9193,-8500,-5291,
-40349,-5676,-1749,-6703,-16501,-17159,-8859,-4566,-11373,-967,-28708,-22515,-6170,4279,-22138,-6713,-15135,-11213,-24576,4937,
-23558,-12640,-12149,-10186,-12832,-20059,-2336,-11921,-13237,-13204,-17014,-20015,-6281,-4223,-18244,-9890,-32370,-6727,-28319,-13155,
-17160,-4406,-20520,-4651,-20665,-19144,-5668,-8628,-4410,-6326,-9083,-13364,-5950,-6873,-27246,-9087,-41748,-17230,-31835,-8044,
-14871,-15176,-13936,-7217,-15333,-22211,-7531,-18098,-10974,-10020,-23245,-19847,-13846,-9752,-9581,-11874,-30448,-10453,-18080,-8823,
3477,489,-14831,-7089,-7141,-17373,-7036,-14446,-4864,-3241,-8047,-8708,-7485,-6823,-25093,-1966,-33904,-10145,-24110,-9994,
21668,2547,-17045,-1838,-7303,-7522,3102,-19166,-1763,-600,1317,-11052,-14859,-11719,-39117,-1928,-26505,-3916,-13023,5379,
38407,10978,-18996,-734,-9925,-15257,12737,-13528,13742,3902,13553,-24445,-10143,-8765,-59246,-1990,-4442,-12630,-3386,5441,
51291,11054,-13746,5054,-3119,-12775,10531,-9915,21966,7403,24286,-22997,-13750,-9628,-83526,-7514,504,-14073,-9101,5339,
63057,14169,-5768,14140,-11113,-10703,-1494,-723,22656,4714,35696,-19451,-8058,-10509,-93263,-9788,-2619,-14432,1301,1807,
33512,9440,-9644,3557,-5075,-4526,-419,-2044,23884,11152,40305,-7391,-5589,-9702,-100856,-11420,-3750,-8714,-1900,4016,
20305,641,3152,-12321,-8011,-11608,5054,7883,20039,5557,23576,825,-1516,-11690,-101452,-4415,-946,-2783,-1124,-957,
1870,-5953,-2157,-10250,-945,-8674,716,6851,12897,6271,2768,555,-2521,-797,-86032,-3822,-2081,-5473,4171,6852,
12832,-7164,19,258,-6217,-68,-8016,7133,1107,3346,-11629,3135,-2382,-2796,-45519,1179,-1639,-3148,-1299,5113,
8521,-307,4866,-2456,352,-4731,-17060,1334,-7951,-1491,-13195,3220,3290,2128,-8926,204,-8033,6437,2711,4628,
4442,4346,4688,10910,8376,-114,-16574,-3284,-14012,-4548,-27914,9250,1251,3450,7202,2056,403,-3757,-6838,1965,
-9302,8958,-1393,-3076,7912,4179,-14716,-6452,-14695,-1760,-27300,12108,6277,6088,23607,10879,-748,-5680,-5964,203,
-10035,5638,3825,2820,12401,4761,-12037,-5042,-18063,-1511,-28135,4563,5711,4040,42494,6090,-5576,-2795,-1625,509,
-4012,-715,-1163,5466,16288,-1452,-2838,-4531,-16709,-4639,-35325,-854,2929,4456,16704,8383,-1718,-4603,-1409,6769,
13719,-4140,2320,-434,11210,-3289,7637,-1958,-8165,4626,-30035,7919,3487,2661,-9796,-5085,-8463,6902,2090,-2550,
18019,-1599,-1479,-16244,8447,3493,17215,423,3730,7242,-29922,-3169,1,288,-43092,-3179,-8621,7565,2592,1132,
19841,4693,4037,-12487,5561,-6346,17991,3110,14426,3412,-31273,-4731,1869,-8526,-74644,-17350,-3419,-547,5473,5590,
22817,4482,-7432,-25676,998,2275,22142,-2059,17711,5818,-19188,-4193,1443,-4067,-72897,-22158,1916,5128,-1447,6372,
21946,989,-4737,-20787,-2061,-1722,30168,765,16543,4739,-5668,-10494,-207,-9582,-63218,-29171,4265,789,-1509,7681,
21283,-1322,753,-9722,-6735,-9090,33142,283,11516,1680,11031,-5818,-17981,-10847,-48166,-22302,9864,-2843,-3102,850,
18531,257,-13361,10492,-13587,-17248,19733,-7215,4481,-3253,26473,-16626,-11728,-2377,-43675,-12890,15651,-4228,-321,-5173,
19720,5236,-8533,18940,-15180,-14207,15310,-10699,-1374,-5074,18097,-15152,-19484,-362,-40728,-3563,19590,-12825,-7168,-12938,
2994,-2744,-3688,20209,-7260,-9970,17480,-8125,-8658,-7258,11523,-23557,-22124,1486,-21518,-12913,7522,-12690,-5072,-5088,
-10967,-5210,-8902,1700,-7857,-18648,8688,-11969,-15623,-4882,3664,-7332,-6885,-3538,-25436,-11905,-2151,-6945,-11058,-1804,
-47619,-7248,-1867,-6525,-13086,-19444,-11730,-11427,-12002,216,-19137,-11336,-10483,31,-22838,-15124,-12517,-10683,-21002,-8153,
-16142,-1992,-14274,-2683,-26172,-20327,-5945,-14631,-7390,-13679,-14246,-11712,-11023,-8112,-27576,-3305,-41930,-8043,-27375,-7719,
-19560,-2953,-19741,-5196,-24196,-23307,-6113,-20639,-5448,-6564,-15278,-12651,-9888,-2708,-24270,-8295,-37685,-16571,-25345,-13505,
-20709,-12918,-16119,-2864,-15687,-28482,-5729,-10301,-4539,-5297,-15622,-11187,-12241,-13524,-20670,-16859,-30094,-9946,-26006,-3015,
-8669,-3687,-5183,-5969,-17951,-20823,543,-10797,-12087,-9895,-24764,-14937,-4785,-6296,-14264,-10543,-21144,-10394,-19946,-2391,
22123,8759,-5702,-13915,-14048,-9486,155,-188,3598,-76,-9776,-23167,-7161,-6247,-31294,-11287,-11572,-9922,-19951,1786,
37651,6791,-14636,3682,-20690,-18002,6138,-10823,15666,6391,8764,-12781,-20232,-6632,-52809,-6349,1230,-14204,-2045,4482,
44130,8979,-9491,3135,-11486,-12201,7557,-143,21371,272,20950,-21213,-22739,-3175,-72613,-10491,-400,-12214,3202,8847,
59150,7382,-17875,1462,-17603,-12832,-1958,-2726,20562,3274,31493,-14082,-9472,-207,-86000,149,5150,-9146,1874,3516,
44892,3348,-6591,-4521,-10310,-8067,1055,2611,23377,6335,30915,-6208,-7872,-7000,-90518,-4660,2171,-9814,254,6999,
23137,-1921,-6126,-4550,-3637,-4223,3447,-1528,21741,3460,6903,-6333,-10887,-3529,-101096,-11587,3836,-1804,809,12207,
18743,-6077,-4232,-8582,189,-7523,-2673,9233,14409,3174,-2871,-1730,-6745,1022,-90930,-12318,-4656,2577,5053,8312,
27712,-8072,4563,1860,4874,-3104,-12125,12561,824,4661,-13359,-325,179,-6762,-48294,245,-4944,-4339,-6892,6657,
18274,-3404,-141,-2476,4783,-7585,-17080,4454,-8949,7596,-14868,523,7092,-1539,-13256,4520,-14346,3565,3367,2960,
10331,1818,1871,2118,7812,-4555,-17484,-2258,-11561,4384,-21255,-1057,11104,2105,6093,2391,-9114,5645,-3493,-3078,
4577,1890,6337,5068,10589,2892,-15787,-4330,-15382,4152,-26004,12787,5222,3157,22559,6145,-6542,-4616,-4613,-601,
-11298,7805,1627,3904,4899,3710,-15318,-1632,-13156,-2118,-24532,7851,14008,773,33604,3181,-4491,-2545,-6268,83,
-1806,2607,3399,2368,5137,78,-2388,3809,-9314,-1530,-28822,3940,6684,4436,8922,3324,-2954,-1906,-4837,-5375,
8212,-3085,-1979,-4605,3330,7790,6566,7309,2111,5082,-28253,-3879,6106,2058,-22648,-1642,-8868,-1477,-3481,2435,
18532,-1038,-5932,-10585,6313,-4470,2808,9266,14137,9253,-29752,-7726,6784,-2517,-64173,-1066,-4775,4176,-601,-2943,
16610,1669,-778,-19882,5593,3300,4763,-2385,19855,10590,-29986,2992,-5080,180,-84308,-8031,701,-2499,-4929,4479,
22421,-1557,-6577,-22727,-1932,-6539,15821,7267,18611,11423,-21052,1614,3745,-10672,-74094,-16836,-224,-6643,5743,4845,
17984,-8481,1588,-23411,3092,-8009,31384,-4492,14571,8010,-11301,-10134,-4646,-6974,-60774,-22473,8111,-2341,999,4915,
10760,-11035,-9535,775,-6205,-5446,35419,-4508,6903,4880,4672,-13878,-10926,-12819,-45655,-23647,11733,-3442,1260,-177,
6636,-7211,-8701,11730,-6472,-9526,24143,-10772,-4952,-119,23176,-11775,-16726,-6524,-32384,-9757,9686,-5541,5498,-3236,
6777,-5289,-14160,22157,-6389,-7505,17007,-10020,-10159,-9096,17673,-25170,-17688,460,-35964,-9705,9373,-6560,3427,-3057,
9290,-2183,-17210,17380,-7659,-16888,13435,-8896,-14434,-9654,5657,-12428,-12664,-2816,-38131,-4539,11307,-9158,-989,-11116,
-10226,-9396,-10339,1901,-11281,-14055,2678,-10198,-22622,-7345,-3118,-8642,-12929,-1520,-25597,-6547,-5739,-6678,-2472,-8070,
-54158,-3390,-4865,-4513,-11592,-13544,-12521,-8759,-20231,-6088,-21942,-18451,-4650,-9688,-27987,-5289,-11147,-12108,-21221,-997,
-35964,-15213,-17206,-2207,-19968,-22950,-5559,-21350,-3163,-9354,-19988,-18896,-8947,-12335,-24253,-13521,-22202,-9181,-26484,-894,
-27647,-13469,-17809,-8729,-17813,-14625,-3145,-35206,-10038,-20546,-14193,-30358,-14329,-7026,-17125,-2875,-33624,-19811,-23489,-7783,
-23580,-14261,-11346,-5230,-20333,-28118,-8411,-22121,-4133,-10655,-13935,-23478,-5729,-12614,-16781,-6086,-30626,-15186,-23237,-5242,
-23840,-1814,-15265,-11152,-32760,-13889,-5680,-3961,-18330,5136,-33205,-16461,-14756,-5092,-9035,-15674,-8083,2176,-25457,-356,
23418,1846,-15548,-9340,-24336,-18024,-3247,5562,3499,6356,-25801,-21665,-13926,-8238,-26959,-8095,-1331,-4881,-13046,-2363,
26916,3975,-14821,2925,-16229,-17965,5882,-375,12985,-855,6934,-20434,-14168,-8784,-38515,-15872,5664,-5088,-9802,9015,
38112,5372,-9641,369,-15315,-15329,3520,-4535,15612,7131,18736,-18545,-23076,617,-54844,-7836,4264,-3878,-1929,787,
47972,3054,-13269,2113,-19455,-7431,2365,3087,17650,8852,26853,-14980,-16564,-9223,-70767,-5145,824,-5373,3796,5408,
43285,1540,-13486,-3408,-10707,-8385,2998,135,20261,6662,19137,-5418,-12982,-806,-75627,-9623,9014,-1612,-1274,2180,
38650,-2379,5094,-8797,-5638,-3687,5649,346,15421,7134,-1348,-3753,-11775,-1981,-83565,-9113,7852,-3859,-3949,-221,
23546,-6562,-6966,-9646,-1736,-449,-886,9405,6289,7789,-5506,-4817,3648,-3261,-64351,-11342,-7161,168,4551,6875,
33585,-9099,6846,2732,-683,-1525,-11317,294,-6019,-104,-16275,4694,-3708,-3139,-27578,-2942,-7335,4432,2310,9170,
23323,-5891,2552,1429,8729,-5257,-17003,1463,-13251,6791,-17491,1916,6084,1163,-5775,1964,-14293,4160,2960,2428,
22362,-2802,-2077,6558,7413,-205,-15503,546,-14051,5994,-27490,6933,3691,2309,5762,6009,-6429,771,-3843,-3267,
11513,1953,-5667,3562,7468,-2153,-13005,8111,-13884,-2042,-28096,-917,5969,2693,24621,6773,-5160,55,-3054,-926,
-20549,5506,4353,7417,10729,-2861,-4264,-6772,-12623,1576,-25560,3473,9129,1983,31803,-3213,-4881,-2464,-1498,3039,
-4844,4861,-3176,-4406,-1743,-191,3084,3630,-1277,607,-24042,808,7198,6563,1279,3862,-2856,996,-380,-4579,
6705,-5443,7142,-3613,-1612,352,-816,-559,12624,2092,-19198,-2671,3246,5408,-31404,-6652,-5505,3421,-6575,5696,
18695,-3887,2777,-10063,-7988,-6784,-13811,12584,22521,3147,-19518,-6189,2601,838,-65527,-713,-5402,3118,1165,-1063,
20867,-1728,-5038,-16545,-7397,1825,-10879,4414,25545,8029,-25555,1988,-10311,-2273,-84604,-2585,-729,2052,4908,3406,
17439,-9007,-3842,-27254,-121,176,8618,7936,19574,12168,-21871,391,-9591,-11038,-70653,-5893,2272,-5922,1073,5852,
17138,-16131,-7020,-24479,-4573,-4337,31000,9133,11483,3165,-16665,-7193,-11503,-19096,-58512,-7404,10623,-5627,4783,2467,
3824,-15975,-2407,-3637,-4060,-1445,34448,-2812,1718,-307,3646,-18893,-18005,-17363,-37649,-19704,6992,2195,9904,-1301,
8841,-7906,-347,15057,-5755,-2960,22792,-10335,-10872,-5316,13580,-16638,-14216,-5320,-28896,-17215,12417,-6048,1803,-12681,
12385,-9379,-5412,9594,-6876,-10905,8171,-18964,-18462,-12590,10583,-15001,-16272,2495,-25514,-4217,12438,-4065,1116,-7370,
7396,-8067,-13079,8187,-12997,-12271,2847,-14004,-23730,-19342,-271,-11314,-4697,-1375,-24534,-1746,11350,-15805,-176,-512,
-10580,-2680,-5319,-2993,-13333,-3350,-6206,-5290,-27036,-15222,-14237,-7723,-3517,-2973,-22084,-12555,430,-11637,-11396,-13338,
-17389,-10247,-13221,-4134,-15419,-13267,-6975,-5881,-21874,-6652,-28059,-13908,-13403,-317,-14597,-57,-8655,-6823,-12533,-8873,
-29511,-7340,-9919,-10914,-15966,-16748,-1372,-21217,-14379,-6069,-12812,-20689,-7767,-10735,-20056,-8429,-29004,-12427,-19793,-2194,
-26599,-9434,-9377,-2595,-10875,-23303,-12762,-28703,-7078,-17893,-8598,-23916,-13132,-11375,-21536,-12440,-42347,-16925,-29415,-6896,
-10895,-12357,-20327,-13504,-11759,-10209,-6196,-14634,-4822,-3173,-25142,-28947,-12564,-11871,-4788,-14188,-30481,-11807,-25539,-3296,
-10426,-5005,-7943,-16446,-35611,-22342,-7826,736,-17753,-153,-24296,-18105,-15299,-9786,-14164,-6196,-10590,796,-18804,9247,
14991,-7163,-14671,-16239,-24181,-24096,-13669,11690,-9174,7653,-30606,-20720,-12010,3301,-12754,-15123,2081,-3482,-14623,-2762,
20498,-1568,-8786,-10040,-18099,-18719,5036,8130,1982,2761,4197,-15628,-23042,3930,-19308,-17355,4165,-767,-9973,-574,
22862,4291,-15360,-2840,-21369,-9248,2611,-2786,8378,5681,13405,-14856,-22393,300,-34942,-9241,6315,-1581,1192,5625,
34092,6100,-6900,1254,-23911,-8729,2250,1403,13599,-2190,13396,-12332,-17114,3481,-46644,-12333,14302,-11326,2547,4490,
30436,3954,-4776,-2521,-10038,-8961,5807,-25,11529,7337,11567,-15362,-9101,-919,-53927,-18248,8502,-4450,2119,1467,
30855,403,-7793,-3497,-1118,-14031,6531,4935,2677,5560,-5972,-4503,-279,3293,-48966,-19100,8806,-6445,2347,-3478,
26691,-3634,-6483,-904,8526,-4783,-2138,10442,-10012,6326,-10627,157,1980,-2895,-25147,-9082,333,-1500,-4439,-2319,
23266,-6822,3539,66,9110,3324,-11173,-146,-19319,2621,-13615,-403,6649,-1589,-2573,-3026,-6976,461,-8123,7433,
28552,-2277,1656,8271,3877,9,-16441,-316,-18392,-2541,-26824,-1848,3136,5999,6563,-1721,-6109,2662,1963,-59,
24445,-741,-2130,2087,7912,-3582,-9781,2986,-16917,1340,-28455,-2849,6998,-329,15259,3775,-5294,1264,-2186,419,
4562,6408,-2140,4185,4203,-132,950,3663,-15629,-2099,-30882,1269,150,-1692,28058,2844,165,-935,-4971,-2734,
-21723,11522,7624,-6083,1804,-6420,9652,-3798,-9353,-2935,-21927,5605,-1186,-3817,28345,5128,222,1894,-6129,874,
-5146,1067,595,-1342,428,-10721,11463,4360,4482,1523,-20245,4059,-4186,3474,-7852,1385,1421,858,-5235,-2393,
-3129,-10934,8477,-2221,-9703,-10185,-10573,8801,20300,2561,-7112,3262,-1090,-844,-31051,-4295,-6255,5677,-4464,4146,
2767,-12728,4257,-3303,-3731,-5390,-24850,-38,27494,11141,-12453,-2126,-6112,1740,-62112,-380,-904,4101,-4389,4875,
11501,-13130,-7294,-11119,-6681,-1249,-20301,9933,27569,15425,-18333,2806,-4156,-6647,-78252,-7349,171,-1032,-683,685,
9211,-25089,-4490,-24957,-2469,-5463,-3163,8532,20196,11234,-24500,-9496,-9930,-7397,-62311,-4194,5158,-9438,12050,3568,
-5637,-30645,-6413,-24176,1561,5081,11904,-1321,7973,9860,-12008,-3216,-15018,-22677,-40094,-12390,5293,-4881,10039,4842,
-523,-15717,-2617,-16212,-1255,458,14054,-5636,-6660,-2739,436,-8215,-9525,-18980,-19718,-15536,11952,-7222,2713,-6618,
11192,-6671,-9492,-5272,-2856,2928,8692,-7307,-20551,-12605,1608,-18932,-16755,-6043,-9547,-11220,11877,-3135,5728,-12374,
9093,-18805,-12668,-1309,-2607,4034,4283,-9917,-29488,-14401,2767,-15137,-7527,645,-6050,-14648,6655,-6528,431,-6093,
9532,-9651,-9204,-5407,-4934,-11042,-5208,-15962,-32955,-9810,-6769,-17004,-4129,4528,-8597,-4374,6035,-8444,-456,-14885,
-21376,-11126,-6920,-14729,-4214,-11344,-5807,-2158,-23101,-12622,-23739,-14077,-4490,-6934,-16970,-14164,-2387,-9115,-3929,-10504,
-22228,-11382,-7194,-16226,-18603,-15917,-9648,-10246,-13468,-10399,-26948,-8999,-7421,-7347,-10976,-6165,-7153,-5056,-19803,-1788,
-28876,-14595,-6252,-13147,-16003,-19882,-5857,-15996,-5817,-12446,-22239,-26034,-16787,-14576,-15976,-12341,-28464,-3459,-23563,-2923,
-19878,-1817,-8076,-6977,-18799,-31267,-5381,-19477,-6035,-4190,-13125,-13444,-7271,-14742,-21854,-3427,-37660,-15748,-25308,-10451,
-19273,-11061,-21560,-10552,-9080,-25191,-8822,-38438,-4031,-19036,-22435,-30949,-16955,-14012,-13647,-5035,-20921,-14271,-19768,-14413,
-31685,4001,-11040,-15002,-28731,-19213,-8146,-6495,-18047,14156,-40955,-23985,-17268,-7040,-17235,-11006,-7221,-3796,-15669,5290,
1279,-13828,-6719,-17313,-40587,-24165,-8397,4559,-9243,4286,-43903,-9145,-7605,-11065,-24353,-11517,12336,1161,-21057,-116,
14745,106,-13037,-12226,-21408,-15547,-8139,6846,-19934,4451,-4434,-8812,-10734,1321,-10552,-20259,9787,-4597,-13463,1528,
15783,7169,-6241,-11117,-21194,-9595,-3419,5276,-11488,-698,7130,-17235,-18697,2810,-2408,-11846,12271,-4052,-10937,3054,
21904,12860,-937,-10133,-18821,-11233,2329,741,-6185,1485,10236,-17529,-22125,574,-13883,-10202,12926,1912,-389,-3024,
16848,13632,-7577,-9038,-8141,-2993,4893,4220,-10206,479,5762,-14286,-6793,938,-16304,-14758,13244,-8041,-1890,2459,
13780,10291,-7057,-5082,-3120,4108,2216,3137,-21663,-614,-6207,-8355,-9481,4333,1205,-11983,6962,-7196,2137,1419,
11246,3497,-5121,-2931,9334,-414,-7733,2880,-30693,5559,-6930,3215,1978,4575,17490,-7871,-533,-6136,-1694,-2191,
24345,-407,3404,5593,8521,-5709,-14641,85,-31205,3343,-17145,8969,52,3253,17676,-681,-1410,-5237,331,-4805,
30917,-1085,2160,-4407,8222,-1918,-8012,7106,-26686,-707,-21384,9021,-3206,1845,17972,8093,-2042,-1135,-5074,-3946,
23306,7891,-2648,-522,3365,-4629,1562,5577,-18475,-393,-26005,-5463,5686,-2996,22648,1108,-164,527,24,-5183,
-12111,15465,1921,-3510,6613,-9488,14854,-629,-12230,-3017,-25552,-3124,-643,-6147,30275,914,3317,-4633,-805,4340,
-20980,12254,715,-9285,-8055,-9634,25000,-6175,-3190,-1210,-19848,1424,2250,-2635,20627,121,4846,-1150,1336,3020,
-15516,-7943,-2250,-8775,-16049,-3806,10680,5223,12021,1579,-6783,7417,-262,4038,-9169,-2632,2222,1137,-9432,3306,
-14109,-20491,3433,3228,-4364,-13824,-18145,12848,25410,6534,-3888,2350,-3652,10423,-32225,-7055,1992,-2423,-8607,1504,
-15518,-22335,185,-8259,-1768,-13911,-31916,2252,30560,12350,-4207,-9223,-1033,8166,-51504,-1702,2286,789,-5659,6346,
-6391,-31378,-5189,-8681,-1597,1300,-29859,6558,25874,11314,-16282,-9243,-6076,-3625,-59644,-4898,4829,-3085,2525,6989,
-5229,-40209,-2485,-25584,-1351,7323,-26179,-2489,15448,11869,-18662,-6447,-10293,-14042,-44775,-3473,9316,-1427,4943,-1244,
-1987,-27938,-401,-36675,6654,1495,-12957,-20,3226,-5942,-20135,-9002,-8977,-15103,-28149,-7245,20774,-8834,2048,-10194,
3250,-10031,-6588,-33987,3203,9533,-8295,-5140,-15419,-9672,-14659,-13427,-15547,-10829,-9637,-11692,14674,-11368,9734,-12647,
11510,-5607,-7477,-33820,3302,10493,-2751,-13767,-30800,-9996,-3069,-10134,-12016,-6615,-466,-8378,7477,-3728,1604,-9839,
17268,-11656,-5859,-17782,881,-237,-8157,-10943,-35092,-12532,-10657,-18079,-5229,-2343,-5112,-15032,6038,-6884,35,-12977,
11056,-17180,-3736,-18289,-2964,-5531,-4687,-11800,-28624,-11468,-17231,-18308,-4250,-3169,-14933,-8475,7526,-4797,-7192,-18659,
-11415,-4907,-4681,-27501,-10748,-13751,-6636,-9978,-28857,-12400,-29188,-4180,-6693,-7115,-632,-7101,-2711,834,-1053,-18118,
-13810,-14478,-8917,-10859,-8109,-17242,-11273,-6578,-11560,661,-22017,-20643,-13679,-10464,-6354,-8801,-12572,-5157,-16565,-11883,
-15542,-7594,-13011,-7495,-17193,-20090,-5392,-24913,-6075,-6776,-10714,-18467,-5692,-5409,-5388,-12579,-26939,-11583,-27949,-13027,
-16161,-14230,-20592,-9114,-13314,-23791,-10119,-52831,-10504,-21774,-18474,-35619,-13486,-17769,-14631,-5498,-34016,-14049,-20110,-17907,
-7372,3004,-18247,-6797,-14248,-17431,5734,-23025,-12775,-6684,-29040,-26316,-14712,-12292,-4055,-8657,-29668,-4531,-15246,-4839,
-20297,-5886,-13288,-10884,-38486,-19821,-6845,2382,-17705,5623,-40422,-13968,-18272,604,-10545,-21007,-6564,771,-11856,6736,
1471,-4831,-4328,-17399,-23056,-21338,-36952,6454,-30892,8442,-41605,-14990,-15868,3895,-4573,-25644,-508,-4091,-9139,4754,
446,6340,-3658,-17920,-25884,-18298,-26750,3807,-39009,1681,-13496,-6791,-16458,-4523,-5873,-12500,10048,-3958,-8720,4258,
6686,14524,-7780,-20823,-18089,-14585,-11843,2790,-36452,6060,2061,-4185,-16318,-152,-5354,-12189,10787,-3282,-8005,1729,
9875,20221,-4863,-5821,-17682,-7604,2854,1421,-37858,8703,-715,-7998,-16290,-6114,-2540,-14269,16308,-5764,-3150,-6504,
4521,19945,-11196,-9258,-7658,-10284,3656,8678,-43240,-2895,7635,-6577,-8643,-5818,18977,-17570,8843,385,3425,4175,
16844,18114,-6947,-5042,-4957,-3509,-57,8652,-44092,-5860,-3178,-8955,-8118,-4199,37288,-11224,5503,3136,6868,-2561,
13254,8373,-9371,-6026,14839,-2184,-7121,514,-40862,5280,-7801,-3102,-1076,6209,33175,-4580,4214,-1964,-2937,-3976,
26152,1336,-8042,-2091,7127,566,-6945,268,-36109,3764,-12618,562,-225,157,27839,2741,1009,4970,625,-4015,
26788,5251,-2297,-3180,4338,-4900,1038,4240,-24948,817,-18705,2697,-5972,2443,25110,1118,378,-2493,6372,-3094,
21062,12648,-6550,400,-3556,-2733,16775,2663,-16223,-470,-26296,-2291,-507,-8220,18615,349,10062,-5544,-3760,-2516,
-12718,17139,-559,-6491,-517,-11241,28415,6093,-8840,4880,-17867,7578,-1589,-11369,26516,-4777,5853,-3717,-884,-6526,
-23033,4026,-1344,-8846,-13645,-9069,29944,-3703,3355,-528,-12956,-96,-247,-3520,13658,-5320,8665,3910,133,2936,
-26710,-22173,-3293,-999,-13219,-13905,5529,12137,15353,2663,-2766,-6076,-6327,10466,-5459,-5420,3065,2592,1531,911,
-25936,-35235,4944,2382,-8865,-10663,-15184,12792,21625,10097,4397,-7033,-1820,7063,-21155,-5747,-2286,-2117,2702,5490,
-15657,-38240,4184,4704,-4734,-9137,-31396,10434,22003,4905,-1249,3254,-9867,268,-33968,-2458,4677,1507,672,3430,
-19569,-40308,1095,-13861,561,-1816,-40680,339,17209,4413,-8729,-15605,-6847,-2222,-34948,3224,6931,1421,5435,1664,
-16608,-28688,-10110,-19900,1245,8794,-43377,743,5827,3429,-19004,-11146,-11315,-15947,-25790,-2410,9559,-1506,10689,-12098,
-11203,-8406,-9715,-38422,10644,10123,-29179,-907,-8017,-4563,-17992,-18978,-3697,-12848,-15052,-12095,10479,-12205,9180,-14208,
5317,1679,-1501,-53811,12710,1063,-19485,-14051,-24674,-10941,-16494,-19107,-9166,-3324,-4384,-8546,9019,-12737,14515,-9582,
12110,1817,-5491,-38969,9721,9807,-9099,-13083,-33611,-13113,-13550,-10548,-8294,-4251,-1400,-15584,4965,-11621,-1163,-2484,
21412,-5607,-6347,-25249,2268,2440,-4738,-15555,-34518,-13998,-23905,-19085,-7332,-12390,-9817,-8837,8708,-3472,-3517,-8995,
2819,-4240,-11653,-18716,-1144,-12569,-4262,-5430,-27411,-17053,-28523,-8586,-3159,-16809,-11944,-9795,5868,-8911,590,-7027,
-20831,-9988,-8523,-24474,-4040,-12984,-2390,-7219,-19770,-16959,-39387,-4686,-14068,-6488,-7396,-15261,826,-4230,-6430,-7784,
-8438,-11724,-15663,-14349,-9013,-4018,-13487,-12950,-22016,88,-23862,-14959,-9533,-15265,-5599,-5236,-14043,-1670,-18421,-3006,
-11498,-1833,-7774,-2883,-22901,-24885,-5294,-9352,-1655,-4893,-6381,-14729,-4300,-10857,-15142,-10345,-32270,-11900,-34595,-10760,
-26469,-4278,-13032,-5588,-11959,-25626,-13630,-25703,-8985,-21934,-24171,-34072,-15007,-11020,-13485,-13967,-31357,-19456,-21932,-9540,
-31807,-6637,-6077,-1134,-18261,-15072,-6907,-17295,-8551,-7433,-27349,-22739,-11722,-8441,-23558,-9961,-21386,-13591,-22641,-10291,
-17592,-5679,-2371,-19747,-24657,-21481,-19237,7734,-18174,14055,-51441,-18517,-20824,-38,-12048,-13283,-4423,-5109,-21120,-291,
-1476,-1029,-12099,-12966,-32282,-21666,-32429,16744,-36814,4125,-51434,-6628,-9989,-6253,-4495,-23412,-764,-4743,-6007,4329,
-418,1313,-6326,-21543,-28449,-13043,-33020,907,-41430,3018,-15276,-7754,-13283,1598,-985,-14177,6327,1060,-7056,7349,
5307,15352,-10066,-17222,-23142,-7607,-13728,6054,-40865,10937,-3619,-6394,-12306,-3755,-3029,-16334,4174,1525,-1429,-2594,
-9067,20852,14,-20573,-9595,-17442,-2666,1304,-41995,7450,2316,-10494,-14763,1330,3451,-13898,6331,-7161,3098,4488,
6562,26715,-13164,-16571,-21381,-15206,-2352,2920,-34639,-290,294,-2062,-6002,-3944,39198,-4084,14626,-9,9468,-4553,
14964,23306,-5709,-8184,-10826,-762,-5393,1571,-33641,3,-3356,2122,-958,-6557,32829,-4246,13745,-9745,-187,-669,
28714,14489,2833,-10885,-7583,1903,-3799,-550,-33209,-1514,-7162,-658,-6768,-2011,27400,1979,10382,-1457,-2411,-5598,
25192,10596,-7420,-9044,2979,-4159,73,6076,-26349,3543,-5563,3962,938,-3935,24973,-4114,2841,4736,2517,-5844,
24510,9935,-433,-549,1744,-354,12246,5477,-19340,-1201,-13919,5948,-6641,-6862,20885,-8228,5731,-5719,172,3825,
10288,18190,-570,-9626,-3856,-10555,21712,8529,-10577,42,-15949,4896,-2072,-8310,17499,575,12508,-7798,-1592,-6015,
-12772,12875,-3199,-12190,-6877,-12855,31331,4842,-2459,-3781,-11657,-37,-2936,-6763,19201,-4405,12767,496,-2019,618,
-29704,-14070,4227,2792,-1693,-12135,24173,1508,6432,3378,-4450,-1871,-5797,462,7875,-12171,11396,-2142,-7893,4524,
-32383,-37639,6295,5798,-10252,-5512,5498,-3538,10374,8897,7870,-4331,-6950,6607,-3885,-4510,4698,2575,-1710,6641,
-31014,-43299,2215,8851,-6287,-11858,-14566,3125,11287,7314,12470,-2448,-7854,7595,-10657,-3900,-233,7387,4873,511,
-32594,-37582,5337,6196,116,-614,-33686,7975,10276,-2886,9717,-5114,-5761,-2955,-13585,-286,942,5123,2130,1034,
-31242,-27140,-176,-8752,9929,362,-45524,-3104,6240,-4010,-3825,-9331,-9664,-3914,-18816,4181,6163,-119,6930,-3781,
-18047,-7418,-6042,-23147,17092,6834,-41438,-1809,-2735,-3005,-15725,-14059,-12582,-10080,-20236,856,6896,-6694,11673,-14829,
5566,10144,-6394,-43959,8018,9572,-38413,-9151,-11604,-13362,-20258,-18651,-6691,-9258,-20381,-4962,10147,-6820,8781,-14235,
19348,7036,-5927,-51554,3385,8477,-26979,-12623,-26176,-12472,-22888,-16032,-3823,-9199,-14017,-5155,5802,-16094,11127,-5992,
22953,-5499,-2581,-46786,4444,9578,-18371,-9864,-31107,-13152,-23365,-18025,-2548,-6001,-9142,-9534,3764,-13930,-130,-5584,
15832,-7779,-1691,-39874,3668,-2192,-13291,-16991,-33417,-15633,-27704,-16669,-12250,-10299,-2756,-5692,1131,-2298,1738,-2570,
-155,-4882,-5892,-30033,-6496,1314,-12776,-12964,-29995,-8532,-30573,-17004,-2826,-7304,-400,-6839,471,-4912,-2925,-17165,
-9871,-6956,-9124,-18304,-4667,-10419,-1664,-7140,-25236,-8679,-34584,-16171,819,-8786,-1286,-8085,-976,-10630,-13119,-12243,
-14787,-8446,-11084,-18897,-10482,-13313,-13194,-11238,-11415,-5639,-27019,-12337,-12006,-13552,-11501,-11076,-11371,-8101,-18552,-3887,
-10465,-11690,-9009,-13162,-6644,-23147,-2849,-29610,-13426,-21644,-15574,-32656,-9632,-9319,-6055,-9051,-35991,-16909,-28486,-10490,
-16540,-6463,-19143,-14887,-23044,-17009,-10133,-38633,-6874,-19359,-15895,-29204,-6660,-16617,-11977,-7478,-37204,-16361,-20110,-19593,
-16225,-7775,-6597,-2488,-24004,-23258,-9594,-13364,-4321,-8126,-6596,-12305,-7348,-3322,-30110,-3017,-28135,-9407,-33857,-5425,
-19913,-799,-4901,-14466,-30814,-23537,-21472,4588,-19271,896,-52525,-13310,-17872,-3562,-17259,-14433,-3959,-6560,-12426,9261,
-6041,-6367,-5757,-15635,-27604,-17860,-19322,6366,-17135,9562,-53839,-6254,-6041,-6666,-18157,-20307,3588,-2145,-19813,2992,
-10140,3266,-3795,-17952,-21488,-17762,-28939,5957,-32973,10042,-24131,-13297,-10251,-9511,-12305,-11088,730,-1512,-4669,5188,
-6699,16459,-4105,-8895,-14317,-11645,-15144,4276,-33685,2308,-12583,-10083,-16125,-3292,-2442,-16709,7574,3151,-5527,1373,
5500,24492,-6814,-15228,-14570,-17966,-6813,6270,-30911,-1743,-10146,-5841,-7606,-3895,17952,-4615,16997,307,-4983,-5024,
4696,26959,-1941,-16053,-12100,-2839,-6757,5960,-27243,7317,-1084,-5341,-13140,-7769,33253,-4706,6007,28,1731,-3985,
8426,27632,-2260,-10352,-13478,-4432,-10601,5017,-21856,-888,-101,-4358,-5747,-3467,31234,-9806,6254,-3913,8871,371,
19250,20953,-1746,-9157,-11070,1469,-3548,4032,-20316,-1506,-1222,-3690,-10381,3475,26551,-9827,5875,1242,8896,-4988,
24552,17638,-4310,-7964,-4945,-1292,3265,8771,-16417,1426,-268,1742,-5157,-4032,18583,-6666,5346,-498,4202,-3665,
19430,18761,-5910,-5991,-319,-6607,11677,12109,-12046,-7286,-4892,234,-5248,-7617,15296,-1178,12855,1648,-1403,-1711,
-537,17772,-3912,-5082,-10124,-1251,21873,9876,-6515,-2875,-6578,-425,-8140,-13168,16444,981,8971,-7153,6078,3798,
-6333,-3844,-5228,-670,-5757,-5620,29368,7129,-4577,3540,-2995,-1666,4749,-3371,9182,-2964,14934,-9133,-5463,-3585,
-31092,-27041,-8676,2571,-6057,-11378,19407,1515,-891,511,10203,-8458,2622,5767,12044,-1579,7918,4035,4531,2840,
-33108,-38864,65,5120,-6409,-4263,4759,12170,-448,-3850,17914,780,-4479,4484,2324,5704,5887,4732,-5595,-3809,
-40531,-37926,-4244,9537,548,-10303,-14461,-514,-989,-3022,18179,7649,-587,3835,-3783,8142,3287,1420,4571,173,
-47720,-25103,3994,5573,14115,5964,-32644,2155,1886,-2681,14983,-1550,-2841,1349,-5719,1778,-1045,-4336,-802,-6445,
-26896,-8815,-7096,-7484,15547,5289,-44609,-7022,1986,-6032,1335,-14934,2251,-7940,-20958,5089,4708,1132,-70,-10582,
-7767,5235,-6497,-23229,13153,8267,-33930,-10379,-1378,-2325,-12943,-8769,-9646,-3702,-28835,-6161,532,-9731,11572,-15012,
17827,3949,-8533,-36326,11943,9221,-36244,-14319,-11500,-7530,-21688,-10944,-2715,-8300,-33497,-3459,6826,-11537,3064,-11362,
21731,7533,-11149,-42155,13609,13248,-25781,-10518,-21883,-6616,-24778,-9841,-6695,-6813,-25340,-11799,-999,-15239,3159,-1056,
29809,1640,-7180,-48611,4937,1788,-10172,-9715,-27520,-14347,-29781,-9249,-3155,-9433,-18719,-6572,1921,-12437,-1546,-755,
12502,923,-3299,-36922,-2165,4880,-1673,-15959,-24456,-6594,-32803,-16983,-6475,-7149,-8713,-16283,-2897,-7532,2356,-9681,
721,-5821,-2664,-24219,-7294,-4262,-8641,-9826,-27944,-11395,-29219,-6091,-8427,-10641,4211,-9814,-3702,-3222,-2535,-15376,
-12633,5010,-9696,-19434,-2760,-12704,-5704,-10496,-23302,-7860,-29481,-6085,-10042,-8789,1576,-9144,-5783,-3025,-13726,-9686,
-4355,-13857,-14443,-7633,-12285,-23475,-7642,-15187,-6472,-4014,-10967,-18016,-5967,-9286,-13319,-4744,-16559,-2612,-24696,-9240,
-20944,-9364,-17447,-15677,-11097,-10134,-418,-35032,-16272,-17751,-12754,-29172,-17594,-10020,-13805,-16821,-33172,-6133,-27680,-5704,
-16672,-8619,-12270,-7694,-21882,-17323,-8888,-20705,-4020,-9441,-20857,-28447,-5858,-18403,-16042,-16780,-36696,-10098,-28414,-19257,
-14001,-15482,-10079,-2349,-16667,-26519,-4029,-19562,-14314,-20184,-17753,-19558,-14312,-16445,-13129,-3161,-34714,-17058,-27120,-9424,
-21470,1721,-2598,-11948,-25277,-14492,-14086,-5725,-16507,9034,-45485,-17303,-16877,-7440,-17942,-15603,-10899,-6579,-18177,9979,
-7097,-4212,-10044,-5564,-37120,-21312,-17910,7082,-10902,3204,-47548,-12801,-5593,-3568,-25215,-9025,8387,-7093,-17796,-4250,
-1942,3843,-13000,-13384,-23751,-20818,-18497,4506,-22652,5876,-30288,-2013,-4741,-11029,-13000,-7559,4675,-3404,-9913,6170,
-13731,7994,-1921,-9975,-12026,-12546,-8015,1483,-34499,9085,-7653,-8540,-6658,-135,-3189,-16246,-1110,-1948,-6973,4610,
7218,18071,-9762,-8538,-10481,-18547,-6434,4894,-27009,10564,-9438,1275,-5469,-6034,22501,-3391,4738,-8560,295,-1315,
6444,22180,-6232,-9998,-5779,-12410,-9771,3833,-22495,1298,-2972,1488,-1826,-3769,25662,-3809,9272,-7353,-8019,3703,
10060,23677,-74,-8100,641,-4634,-8317,263,-22072,5411,3375,1311,-10641,-8314,25476,-3971,2042,3512,-4542,1905,
18259,24890,3799,-12904,2963,-3424,-4997,12830,-18835,32,6908,596,-10834,502,20263,-1410,2691,-193,-5365,-7535,
23770,25002,-4334,-9923,-1169,-7328,792,9746,-18118,1905,8470,3564,4569,-9093,14014,7771,6223,-3053,-2938,-7665,
15013,22304,-2185,-769,-7565,-4129,7216,6914,-15003,-2857,7942,4460,3791,-10130,15051,5695,6501,-5103,3373,-4921,
645,13116,-7457,10849,3140,-5628,15011,5079,-11003,946,6467,10795,-4369,-17397,10224,-492,5758,-1995,-1586,434,
-9848,-8601,-2777,4786,-2627,-10197,18614,2080,-10371,2177,10257,3751,-1830,-4995,10338,9671,5124,-6626,3835,-2040,
-31276,-26056,-226,9203,3156,-6290,11802,282,-7455,-7036,20162,4628,4560,5550,11489,-2961,4729,-674,-5538,3033,
-39462,-35834,-4486,11177,867,164,2268,-3873,-9491,-4257,21881,-4094,-162,7408,7296,7890,-934,6025,2433,-3434,
-44822,-28592,1244,11352,9081,-7439,-15680,-5043,-3761,-8237,21533,4214,1142,2514,-1394,4949,-2501,3870,5110,-6383,
-35694,-15217,5757,6011,11873,-839,-32011,-4685,4058,-11906,8490,-5475,-5250,6542,-11139,4424,818,-4068,4766,-15071,
-16978,924,1984,-731,11285,-287,-40900,-9270,4180,-6684,1278,-3431,-10043,-10411,-24710,749,-5927,-3205,9269,-13809,
1290,8918,-2577,-16992,16886,6320,-43021,-18704,268,-8700,-10496,-12920,-2283,-7968,-37496,-4578,-1657,-12193,159,-1110,
20393,-347,-10427,-30841,9850,9739,-21689,-18217,-6868,-4731,-21603,-14740,-9715,-9119,-40707,-6055,-7150,-7759,9953,269,
26572,-222,-15382,-25020,8151,7269,-12993,-26179,-11154,-911,-33920,-20690,-9216,-4745,-35415,-18053,-3776,-5650,7697,1549,
25087,184,-4196,-26124,3191,2588,-4649,-18771,-17614,-5073,-35134,-14699,-2262,-10335,-23419,-15333,-2447,-17267,641,1018,
14642,3367,-6774,-27665,-3478,-4858,-2068,-8447,-23167,-8137,-23754,-8571,-692,-15562,-10396,-5749,-8805,-15187,879,-2619,
-6504,-8084,-8624,-23681,-3161,-8115,-4950,-10283,-14963,-2786,-20201,-8508,-6203,-8103,-9172,-17208,-8187,-10720,-6641,-9360,
-6739,-6645,-14280,-6794,-8065,-22684,-11506,-13887,-9512,-8930,-11805,-20905,-7173,-10094,-9132,-5519,-9463,-1246,-10891,-3041,
1925,-15851,-14418,-5408,-11100,-20448,-3370,-16534,-10090,-10025,-11134,-13492,-5593,-9008,-10726,-6456,-26574,-13347,-30039,-4275,
-29284,-4069,-16926,-15357,-22503,-11951,-9707,-19286,-9213,-13579,-5238,-22502,-16811,-8727,-17196,-10082,-36458,-13107,-25581,-8219,
-26988,-5945,-16192,-15005,-20214,-16192,-13567,-24475,-2185,-6226,-20252,-12395,-17618,-7302,-19865,-9002,-33448,-5452,-33801,-11931,
-22177,-11212,-21910,-5119,-17252,-16892,-6595,-39247,-7331,-23328,-21429,-32808,-17513,-13089,-19549,-14914,-31138,-14015,-19943,-15710,
-27989,513,-14455,-4566,-28991,-14379,-10632,-5977,-18390,3551,-37632,-23393,-9052,1901,-22714,-6239,-14332,-9604,-15621,597,
-9766,959,-1653,-15149,-26512,-27401,-15508,558,-14687,5758,-34425,-14329,-17052,81,-19645,-2954,-4865,-4221,-18593,-683,
-5205,2215,-2094,-7016,-17769,-25090,-7788,9618,-27491,5998,-23319,-5557,-11645,-7044,-18696,-6925,-5660,-6541,-14715,3892,
509,12074,-8355,456,-19730,-18216,-7049,4,-23422,3666,-17779,-2030,-5585,-9042,-10387,-6055,3043,-6478,-12698,6878,
11275,15489,-8492,-10344,-4352,-20737,-7490,6948,-23553,10378,-3044,-3748,-10587,2980,15799,-675,-4566,-4986,-3156,-1011,
10484,18015,-7805,-9446,-8395,-9437,-5861,4217,-22326,4522,4440,-6167,-4921,-824,22944,-2415,-4597,4465,-3272,1011,
18093,20445,2148,-1338,1412,-11974,-5578,3098,-19256,9922,5826,702,-6950,-3792,16633,-5339,-4014,741,-4234,-4870,
20503,21014,-1140,1689,4448,-11439,-3486,12246,-17346,3900,6633,-598,-9886,-6046,13025,-912,-5548,-5027,-1294,904,
17206,20434,-3861,855,193,1718,-745,5813,-15282,790,10901,918,2402,-6508,10428,2632,-1035,-4783,-6626,2996,
17269,15509,-7031,11799,-3340,-8577,5258,3480,-14477,-3047,6093,9669,-3171,-16282,5536,10615,3243,-3756,-587,2540,
2560,3531,881,9348,3467,-6677,12385,5882,-11623,-2478,12346,10490,-920,-14967,5987,3146,-2451,-3185,-681,3408,
-5149,-9530,-7256,5897,2696,-8389,10367,7041,-8152,-12976,15154,5391,10706,-2709,1090,3296,5083,-1684,-10963,2303,
-18268,-27242,2116,12784,3073,-8488,9426,-2339,-10858,-8010,17248,6875,2201,6747,4365,3544,-500,-887,-771,-5714,
-35390,-35085,3518,16759,11463,-2125,843,3189,-8751,-5311,22140,7387,-2991,4995,-1330,1295,-7648,-3736,-5919,-9939,
-44008,-30471,-3291,10676,8401,5359,-15379,-4694,-793,-10154,20543,3150,325,851,-10332,6884,-9478,-3388,404,-3196,
-33778,-21942,-795,11119,10566,8477,-30837,-8988,5681,-7798,13183,-9274,1737,-1365,-21114,1194,-10294,-7483,-2175,-10893,
-6951,-7478,-11451,-2513,14447,-3511,-45557,-15937,5445,-12240,5396,-13441,4358,-2324,-38331,1683,-11922,-641,3755,-10941,
9368,-15968,-11132,-14584,16822,12304,-43558,-21415,3498,-5456,-9493,-7944,-7719,-4031,-52625,-3542,-14535,-8564,-1128,-4751,
27646,-11004,-6407,-17445,6995,-335,-28385,-30584,-4516,-1268,-22408,-11341,-3788,-13173,-49058,-4812,-15858,-13593,7995,1670,
36327,-4481,-7123,-22829,7665,5776,-7768,-20086,-9642,-1375,-28941,-14409,-6898,-5326,-44243,-9128,-11156,-15549,-4023,-3075,
27966,3,-6582,-13302,6893,-3005,1783,-15394,-11119,-1480,-21463,-5817,-10604,-13338,-32956,-17519,-14624,-12396,-4379,-1562,
15006,-703,-12106,-21374,-941,-7746,-1378,-17066,-12298,-6175,-17499,-16449,-9620,-8413,-21905,-3958,-15069,-14238,1291,-370,
10466,4402,-2896,-13721,-13370,-13001,2669,-22853,-8608,-3474,-12929,-19973,-7674,-2866,-7234,-14552,-12300,-10933,-7333,-8846,
-6981,-5816,-16254,-3295,-7494,-8979,-3194,-19426,-12490,-6212,-13370,-18097,-5994,-8028,-8121,-10220,-24432,-12570,-19005,-10567,
-11656,-6601,-12209,-13872,-8009,-11613,-11357,-20213,-2063,-6793,-16558,-26694,-17771,-6974,-6198,-8971,-35814,-17283,-27265,-7207,
-20826,-13300,-10565,-7357,-24495,-21008,-117,-19300,-5741,-4393,-8352,-18074,-8946,-14490,-23770,-5705,-38443,-16769,-32168,-5206,
-24346,-5557,-15583,-4129,-22972,-16105,-10878,-42199,-13713,-26287,-25119,-30736,-6254,-16463,-19172,-6830,-35965,-19939,-19196,-19620,
-25852,-7789,-17720,-12776,-18237,-22078,-13984,-31745,-9522,-21258,-21033,-31913,-12052,-13440,-16118,-5499,-39059,-11756,-18521,-11777,
-39284,-2419,-18618,-12477,-13733,-10336,-7763,-12786,-7319,-2152,-29001,-28453,-12294,-11976,-16847,-12409,-20487,-12717,-25177,-324,
-16223,10298,-5805,-838,-29238,-26626,-7050,-1340,-14842,-2310,-37158,-17172,-4111,-2647,-19737,-14588,-10671,-27,-19836,-4661,
-5620,5215,-6705,-3080,-22260,-26668,1446,1477,-21917,8989,-20040,-10809,-5037,-64,-21425,-8860,-9032,-8022,-18821,1392,
1178,10816,-5107,4964,-15879,-14627,208,3818,-25641,8134,-15539,-4066,-12961,-3179,-11248,-10914,-11024,-5556,-17609,3739,
26171,12738,-5650,2630,-8982,-20379,2122,8595,-25631,-318,-5768,-7494,-6513,-6152,3430,-5518,-8877,-2000,-14463,7879,
23277,16838,-4592,1834,-9902,-17135,-1337,5924,-21801,209,2986,-3579,-8908,-4690,9176,-500,-8734,989,-12974,4123,
22086,20006,-7970,9384,-8294,-6021,-2376,1872,-19558,4648,6589,-2822,-7674,-6775,7663,-1283,-10623,3074,-8532,2748,
17249,19363,-13729,337,-7094,-5929,2192,6792,-17999,113,13941,6279,3544,-3884,8667,-3450,-11926,1068,-9280,4920,
21082,18950,-1176,3736,-10753,-8870,246,994,-12794,-4485,11619,7802,-3040,-1299,1703,5194,-6689,-1316,-5177,430,
18788,7716,539,-11,-4816,-13589,7733,10069,-10560,-5702,14142,11173,4509,-5781,-4950,6957,-7000,-7146,-8832,2504,
8908,-4257,-8124,6991,6506,-3196,6715,2802,-5485,3325,12330,-573,-1021,3551,-12828,3495,-6842,-2218,-12762,-208,
6441,-15754,-706,12757,4073,-11597,4731,2617,-2903,-4658,12681,3965,-2781,-773,-16906,6826,-5095,-2089,-9760,234,
-7327,-32566,-671,12952,544,921,5027,5069,-26,-11228,16353,-3080,-6164,7084,-15361,-1160,-14466,-2214,-515,7458,
-17564,-47257,-2292,13982,11230,-9396,2320,-3554,-121,-4022,19647,-4664,-4526,-426,-25899,5457,-16874,68,-2929,2587,
-22713,-47743,-2984,4433,5262,-3247,-13165,-4059,9080,-13796,23317,-3141,2249,3366,-34411,-1197,-18868,2128,-4786,-2172,
-16943,-38885,-4437,4053,5340,5007,-31209,-9878,3867,-16773,23972,-567,2112,3272,-43835,5566,-29606,-3547,-1515,-12056,
-6266,-21057,-5896,2802,8235,8455,-43924,-22020,5687,-18537,12038,2866,-2707,-5562,-64585,2963,-34752,-10774,-351,-13096,
15712,-18121,-14124,565,8054,5122,-35003,-37439,2752,-26036,-8174,-3623,1285,-9606,-72111,4429,-28787,-15875,-1597,-18795,
29003,-12074,-3283,-8459,8175,1910,-20152,-42031,4489,-20741,-15081,-15466,-4203,-12202,-70335,-792,-25562,-20568,-2678,-6038,
34623,-1198,-9717,-8429,-1670,3519,-3093,-42367,836,-10441,-15781,-9107,-4915,-13597,-56844,-10142,-21108,-21024,-2461,-5861,
29309,-3646,-19778,-12271,-3287,2565,-2595,-22931,-1107,-10426,-4673,-19816,-2112,-7962,-46445,-7118,-19293,-22295,-10259,-4176,
16206,5417,-8263,-14449,1567,-11810,2456,-28471,-5078,-10596,-4639,-14287,-7737,-10511,-25722,-5997,-19444,-20160,-13335,-3132,
10467,423,-10063,-9378,-7393,-9559,-8566,-14328,-8450,-13357,10059,-19966,-3378,-7557,-21647,-9083,-30762,-4636,-19785,-9235,
-10329,-8024,-18610,-7517,-19490,-13094,259,-18281,-2781,-11632,-8455,-21228,-4347,-12772,-21977,-5490,-30794,-1959,-26062,-12989,
-26844,-11642,-10044,-14900,-18529,-25266,-12294,-14731,-6829,-6260,-17492,-18132,-9108,-10864,-12366,-11947,-32735,-8332,-29988,-7004,
-20923,-9200,-15938,-14800,-16475,-13843,-5209,-18034,-12182,-8258,-15978,-15886,-14119,-15675,-13591,-10249,-38100,-7101,-33425,-5210,
-26038,-13710,-20494,-7443,-15577,-29969,-13022,-22163,-4528,-12443,-12534,-22239,-6658,-5475,-19199,-12022,-40376,-8351,-24982,-5297,
-21961,-14498,-13731,-3924,-22962,-23539,-9694,-14291,-4551,-6811,-12289,-13566,-12576,-5715,-17561,-15682,-38875,-8359,-31000,-4250,
-14435,-7547,-11888,-6038,-22828,-21519,-4074,-13125,-4317,-3816,-8812,-22251,-14890,-3108,-24432,-4983,-42147,-12228,-25852,-9828,
-19136,-10068,-7884,-12889,-15869,-15934,-121,-5110,-10249,-13308,-25935,-16369,-16187,-2196,-17148,-7782,-28642,-3788,-26861,346,
-9817,24090,-3011,-2472,-25502,-20410,2089,-12620,-27664,726,-31196,-12058,-13008,2103,-19087,-2561,-17523,-6383,-21398,5482,
-3002,14855,-4672,-5405,-32525,-26988,1397,-91,-23949,7500,-20056,-3836,-5724,1923,-28352,-1975,-15712,-8852,-34939,6506,
6151,20342,-11329,2991,-26850,-22066,2171,6568,-26266,4426,-6464,626,-15884,6787,-26180,-6892,-21637,-5603,-19968,4765,
16911,19544,711,-5384,-33132,-32361,-4068,10530,-15406,11784,252,-11082,-870,4335,-19550,-7226,-27643,-1348,-19940,-1648,
22791,17760,-7479,8973,-21249,-19186,3831,13765,-16925,3869,5920,-4586,-1660,-544,-16285,-11976,-23866,-2837,-22339,4657,
23478,20059,-2833,-4448,-24751,-22353,8086,5998,-14471,5806,16454,2669,1173,-5818,-6675,1963,-27363,-2482,-14169,1539,
11375,13687,-10800,2166,-17708,-20116,4560,6291,-4048,7834,20280,384,2334,-4222,-13037,195,-29012,-2406,-11715,5369,
8988,2615,-1745,671,-9091,-23158,12330,10507,-2161,-1713,18954,706,2873,275,-19683,-5146,-27620,-147,-16760,1122,
-2016,-3536,-11050,1217,-8914,-11059,5170,-1262,7449,-1550,14247,-7547,3299,5870,-33681,484,-24691,2210,-16756,5312,
-6027,-21614,-9021,7257,-8873,-14600,5443,3560,6879,4604,13390,2599,2854,-5659,-38158,4903,-32444,1109,-15605,1778,
-11013,-43363,-6951,2106,-2485,-7744,7329,10880,7274,114,11553,-3676,2494,-3801,-42696,3789,-44900,-1034,-11420,11631,
-12398,-52808,-585,1588,-1595,-10202,2087,-1704,4305,-7737,-1093,-3953,256,6313,-57801,1723,-52275,3964,-8419,-1980,
-38093,-39050,1304,-650,12810,2207,-10084,-9268,4193,-6151,-5437,-7446,482,4533,-63088,-2875,-67910,666,-2440,-4225,
-16092,-35696,-6328,1966,-1576,5177,-23012,-10273,8249,-22876,-18041,1262,-54,1412,-78310,785,-61954,-6503,3204,-13770,
-6138,-22380,-5663,5816,13098,-5723,-32440,-25616,4957,-22010,-15932,-4497,6116,-5520,-81557,-1258,-60147,-10850,-597,-21420,
9816,-10647,-15288,5166,14570,3162,-26977,-39636,6828,-35813,-18429,-1077,-3328,-7015,-76434,-5554,-45856,-9121,-9589,-26237,
22384,-10816,-6336,-8351,7500,3350,-6839,-43796,5871,-17714,-10114,-5458,-7515,-13547,-68583,-4924,-40685,-14660,-9547,-20165,
20927,4982,-19135,-5570,1584,1650,-326,-51135,-363,-19609,-8978,-6149,-7066,-12411,-51164,-6590,-31929,-22157,-3834,-13413,
20608,1038,-19424,-12028,-6112,-2175,-5908,-37704,1005,-14549,1365,-20983,-4768,-4025,-44392,-5130,-27003,-21881,-11004,-4854,
16353,-10864,-13744,-10325,-3250,-12205,-9968,-32943,-7566,-4021,-1144,-22840,-10019,-4496,-28240,-6048,-26444,-12527,-13046,-11324,
-1565,2660,-16035,-3492,-13797,-21793,1798,-20010,-3095,-11636,-6172,-15014,-5417,-9170,-24830,-11023,-26535,-17696,-16168,-6829,
-21385,-8148,-17562,-12297,-20144,-19613,-9271,-22163,-9345,-9762,-12292,-22093,-12024,-16611,-13014,-6959,-36188,-6019,-23068,-5607,
-28420,-9444,-16264,-8504,-20832,-24161,780,-35338,-13280,-19238,-28276,-32334,-3938,-17605,-16546,-7670,-29051,-20560,-17263,-16491,
-16999,-3639,-12571,-5608,-22266,-17891,-4377,-12954,-9309,-15585,-9645,-21426,-5376,-4314,-21102,-8468,-43289,-12802,-33632,-2628,
-17138,-12163,-17078,-5830,-22387,-28619,-1431,-10043,-4055,-8441,-16387,-21640,-7664,-8593,-23929,-5349,-39279,-9718,-34554,-12811,
-18029,-6037,-9902,-5743,-25582,-29649,-11362,-16722,-11531,-17824,-13245,-15410,-4090,-3940,-13129,-16430,-34219,-6286,-28927,-4635,
-27977,-18040,-20577,-11303,-13991,-18749,-3537,-40889,-11918,-17394,-23002,-28294,-13681,-14866,-11967,-17131,-30389,-21925,-21372,-8627,
-18288,-1390,-17482,-6658,-18672,-22475,-5987,-20855,-7773,-17961,-15299,-22496,-13494,-6648,-22033,-7029,-42761,-14370,-21861,-9762,
-28580,7011,-13311,4647,-31726,-23135,2291,-11547,-13131,3539,-30225,-14973,-5138,-4513,-28495,-3713,-23334,-81,-24499,2382,
-18945,17049,-2498,3346,-41884,-37018,-4872,8088,-11992,3490,-16927,-16007,-16089,2311,-33251,-5434,-24970,-4487,-28030,1638,
-15521,5527,-4903,-7105,-55538,-39478,8293,11703,-17754,4337,-23045,-7138,-5157,2422,-40331,-2142,-20504,-3919,-42029,5692,
-3257,20383,-12103,5049,-48710,-36390,1058,5880,-17747,14436,-8516,-7081,-10194,-2947,-37571,-2715,-30789,-7230,-39958,10888,
-4141,16886,-11064,6125,-57712,-29575,1696,1255,-20717,10918,1304,-6760,-5462,2016,-38056,-1616,-39498,3202,-38600,6393,
-5812,22880,-7371,6282,-42654,-24663,4538,5155,-10070,6762,-8996,-9427,-9980,4415,-30611,-3042,-43433,-6703,-26596,1966,
2357,13917,-7828,4851,-32380,-26340,4218,6741,-2297,-1813,6062,-1160,-1094,-726,-24408,-3436,-52890,2896,-28874,2619,
-16221,7485,-12128,5752,-22185,-12855,19148,1534,7709,-5726,-1190,-5580,136,-2494,-38960,-4640,-48399,-11344,-27506,6319,
-25003,-2988,-3791,7153,-13611,-21447,16175,-9144,6107,-10098,-15130,2761,2351,-1853,-44997,-1523,-65136,-1720,-27161,-869,
-32350,-16809,-9806,15908,-13529,-10869,11180,-3117,10824,-11228,-6689,-1844,-5267,-2759,-53543,-953,-71628,2525,-24079,-4646,
-38339,-32628,-9415,16770,-3159,-12950,12805,-13371,4595,-10605,-9588,-309,-2220,98,-59018,-1323,-75779,1726,-18133,-221,
-47610,-40862,-10970,3583,-2721,-12080,11214,184,3254,-18622,-18703,-268,4993,1681,-59607,-1799,-82888,-5459,-8979,-2778,
-40548,-48431,1132,640,3623,-10776,-1948,-1416,4015,-22762,-20163,-820,-2016,-4864,-65262,5546,-77780,-6577,-12427,-10542,
-34219,-33868,-5924,556,982,-8281,-13296,-13476,9459,-29713,-17565,-1323,-2086,-6577,-63613,-2473,-70656,-1440,-4211,-10838,
-10805,-15382,-8011,-7567,10025,-7995,-18279,-19890,8101,-12910,-15036,-13278,-2042,-5505,-57482,-1132,-62760,-3616,-6766,-15733,
7861,-5021,-15448,1820,1364,-6696,-21647,-34002,6422,-31526,-18208,-9712,-438,-4946,-56728,-1750,-43898,-17262,-8901,-22766,
13348,-16083,-12664,-4253,1666,-10167,-11110,-47939,3987,-22830,-14647,-14877,-2872,-7179,-48843,-9990,-37959,-21258,-2960,-12499,
12601,-4704,-20263,-12688,-1400,-12777,-3418,-30719,1661,-10596,-4782,-20177,-5533,-11432,-37262,-6354,-30331,-17470,-10605,-10571,
8802,-2413,-8801,-5671,-1441,-12041,2622,-35451,-7681,-14098,-928,-24832,-8110,-11043,-24932,-14384,-31437,-8422,-16262,-9199,
-13528,-2879,-17352,-13767,-12049,-12903,-4086,-33182,-10818,-16824,-14045,-28633,-6041,-5964,-15508,-6240,-28625,-15016,-20204,-12344,
-13192,-9428,-10555,-4224,-23087,-16704,-12478,-24357,-14659,-18001,-18339,-27805,-10342,-3924,-15704,-10620,-35669,-11049,-26483,-18927,
-17485,-6109,-13443,-3420,-22495,-23067,-6289,-23400,-11551,-9589,-11644,-17899,-17259,-12689,-16781,-6716,-39570,-13729,-19763,-15822,
-25999,-17598,-15148,-15755,-19327,-14376,-11793,-39565,-11937,-14039,-19763,-35549,-12415,-14751,-14753,-5122,-33099,-13052,-23650,-16930,
-17943,-17385,-13045,-4243,-18504,-20427,-3190,-23259,-12224,-21438,-15755,-29977,-12305,-8453,-19576,-7699,-42897,-20589,-19954,-15485,
-26200,-6097,-10457,-11011,-19515,-17302,-6788,-30862,-16089,-12907,-19774,-18951,-19234,-6654,-7444,-14384,-35625,-14709,-20786,-8512,
-20176,-10043,-22437,-11329,-22623,-25292,-7994,-23608,-8955,-11681,-18792,-24210,-5279,-10624,-15368,-11313,-33173,-10660,-25681,-9015,
-24161,-10144,-19752,-12763,-18881,-24049,-4149,-18909,-5633,-8746,-18601,-14287,-11544,-14603,-17432,-6830,-34411,-10195,-30971,-10561,
-21304,-1799,-16516,-6120,-12569,-28926,-5162,-12363,-10712,-7521,-11891,-9248,-12470,-6426,-13503,-15421,-41990,-9595,-31214,-3259,
-29616,-10479,-15258,-2621,-16982,-21729,-8211,-26903,-9259,-4874,-15895,-21359,-14708,-8618,-13324,-8729,-32047,-15629,-21121,-2663,
-26728,-3459,-16596,2625,-20421,-19197,5489,-8820,-8167,-7889,-18181,-24237,-3033,-5132,-22498,-4874,-36481,-9451,-24725,-4478,
-23441,16063,-10601,-4355,-31134,-22589,8074,-5867,-13044,1647,-13288,-11178,-7894,-682,-22340,-5677,-43287,-7517,-30014,4587,
-21610,3962,-1618,-3726,-36803,-29056,5741,-4682,-3804,84,-7653,-10357,-3936,-4478,-44043,-2446,-41008,907,-42743,-343,
-21065,21323,-9272,5790,-39587,-27974,6464,-7447,-7327,740,-21542,-17470,-12207,2855,-33841,-5298,-45963,-7815,-26348,502,
-17484,19652,-9509,-2505,-22178,-23165,10719,-5297,-7519,-2502,-13381,-16666,-15367,-1374,-28244,-2641,-67999,-5063,-28410,8435,
-16757,15118,-7282,3159,-19451,-26771,13103,-9687,-2090,-8809,-15407,-4471,-8088,-443,-35312,-6288,-62942,-9093,-32941,7099,
-21541,5383,-7930,8499,-25791,-20438,14713,-7386,755,-7376,-15312,-6408,-12801,-8218,-34656,-1960,-75656,-514,-35990,-836,
-22512,5763,-7993,11835,-17982,-12668,7857,-8093,-1849,-15921,-17785,-13680,-8107,5784,-30948,-8006,-81762,-4314,-22585,1069,
-37750,-6602,-3754,-3019,-6563,-11681,13524,-7372,-4689,-5068,-20501,-12071,-891,1004,-36772,2186,-81189,-4095,-30286,-6469,
-39618,-16239,-11708,10066,-9486,-18134,5037,-8098,1817,-3385,-22920,675,108,538,-48690,-8519,-73049,-3726,-22034,-7176,
-49405,-12881,-13035,-3215,-4311,-13083,-374,-4504,2956,-7621,-23580,-12,-1320,3753,-43492,-8061,-80470,-458,-16001,-9208,
-40015,-20189,-1435,-2379,-3584,-15193,3658,-13012,5947,-17202,-36873,-7573,-10057,-1158,-49742,-2516,-66477,-10119,-11485,-13776,
-27048,-20470,-8647,10939,-9422,-9861,-2780,-31679,113,-26033,-43735,-1425,-8356,-5515,-38812,-6605,-57519,-11828,-4117,-16365,
-21836,-12344,-14938,2595,-5863,-958,-7004,-25646,-1147,-26976,-28379,-14575,-5155,-8140,-28730,-7076,-51971,-10032,-8232,-13488,
-4690,-7696,-8398,-4734,-11152,-13559,-8799,-33442,784,-16823,-8587,-6076,-874,-12832,-28385,-7975,-36111,-16149,-17549,-9388,
-5655,-6107,-11776,-9427,-8849,-12715,-5499,-49237,-9089,-34639,-18320,-22709,-10310,-13144,-13376,-8710,-31025,-19227,-8083,-22937,
2153,-7238,-11484,-4214,-17109,-12872,-10103,-18729,-10058,-11849,-3854,-12553,-7197,-14004,-20822,-5666,-34438,-6170,-29027,-3632,
-826,-13653,-14463,-7392,-3676,-20742,-6030,-33496,-15781,-13335,-5333,-25987,-14139,-8287,-10197,-13070,-27522,-20513,-14937,-16551,
-16713,-17530,-23496,-5623,-19119,-17428,-12939,-38802,-4000,-21641,-16010,-32531,-7257,-15398,-23283,-16785,-32553,-18168,-19552,-18842,
-25642,-16368,-13309,-13553,-10617,-28136,-11144,-25513,-6947,-12677,-15622,-15173,-5235,-14745,-19919,-3605,-35154,-17134,-34963,-7287,
-24792,-15821,-11682,-10721,-14734,-24159,-4591,-30289,-10703,-14630,-11452,-23553,-15525,-4736,-16372,-9205,-40333,-7514,-24164,-12438,
-20063,-3089,-19263,-14103,-19160,-19037,-1441,-20250,-9571,-12334,-18497,-16651,-15481,-7483,-19510,-11179,-41645,-11148,-27676,-4484,
-25649,-13865,-14268,-9330,-17846,-22853,-9345,-37041,-15588,-12572,-14270,-21764,-12790,-4393,-12169,-7420,-33450,-18612,-23984,-16445
};
localparam signed [35:0]b[0:783] = {
-11743,-4156,-13228,-4434,-12454,-10903,-7629,-10582,-2338,-7472,-16910,-8392,-2859,-10542,-11685,-13026,-12720,-5187,-8639,-9965,-12557,-2583,-5600,-724,-3658,-16821,-13293,-6774,-3005,-12366,-9426,-6973,-4374,-11477,-12745,-1143,-12445,-12497,-13434,-13156,-12523,-8997,-2336,-8016,-15238,-15227,-7128,-6573,-8337,-5718,-7755,-6100,-3917,-10747,-12818,-4553,-9711,-2501,-6980,-14552,-6883,-5663,-14525,-7119,-12020,2509,-6788,-9803,-5309,475,-10010,-10677,-9938,-15680,-9086,-7661,-7582,-5883,-4047,-3801,-9617,-9499,-13608,-10294,-12227,-11393,-14249,-13841,-6886,-6446,-3013,-4445,401,-6932,-10038,-7491,-7845,-1968,-8384,-13118,-6490,-10083,-15690,-3945,-13854,-17331,-11311,-11558,-14021,-12199,-10262,-13999,-9291,-14616,-11536,-3432,-3717,-11879,-3631,2408,2237,-4521,867,1780,-3009,-3836,3266,-892,-2396,-14882,-2224,-16353,-13673,-12414,-17944,-9256,-7240,-7217,-9239,-16690,-13923,-12898,-1514,-2303,-2878,-1176,4873,2925,3105,367,4654,5996,1650,-5412,-307,-100,-593,-6616,-5596,-5313,-7560,-14363,-2768,-14154,-7171,-4855,-13248,-14030,-5373,-16133,-5715,-631,-2341,-4785,-7190,3967,3159,-169,-2525,3635,-1308,-5857,-8240,2313,-12180,-9709,-1375,-6785,-13724,-5942,-12684,-7039,-10505,-2477,-9584,-14952,-8099,-11281,-3126,-7805,-3059,-7306,4087,3591,3003,-2845,-1867,4091,-842,-5959,-3738,-2245,-10326,-4364,-7560,-7331,-10732,-12469,-18128,-8945,-2226,-2898,-1950,-13043,-9531,-499,-2543,-10710,-4952,-7247,-2281,8695,1986,-3161,-5649,1644,-12054,-15319,-7524,-12202,-6291,-5553,-1544,-8442,-3126,-9293,-13513,-4837,-3142,-5307,-6199,-3933,-5340,-11860,-2866,-1422,-7064,-8405,-5292,2698,3214,2771,-2149,-3444,-15052,-16373,-13571,-12300,1770,-1416,1589,-5167,-7930,-12382,-8526,-9396,-5066,-9761,-15569,-4257,-15302,-8160,-11885,-8883,-9697,1667,-223,-2294,-1723,3858,-6746,-10485,-12530,-8422,-5632,-9104,-1415,-8094,-5506,-31,-17878,-14450,-11153,-11552,-13660,-11649,-17667,-14822,-12702,-2275,-2796,489,-7834,-3929,-9362,-9562,2365,-7025,-3291,-12155,-11337,-8109,-9220,1772,-5951,4621,2827,4618,-6850,-15108,-17893,-11332,-18530,-14658,-6177,-14457,-13092,-6040,-3751,-3144,-6429,-11983,-4519,-7186,-513,-7347,-9592,195,-6830,-4948,-9116,1337,6275,4198,0,-2444,-4731,-8100,-8999,-7921,-12652,-10284,-7949,-12577,-8440,-5890,-12920,1161,-8092,-13736,-6197,-4797,-994,-4020,-2620,-3306,-4298,5917,-4606,4765,3773,-177,7736,-1252,-5806,-6984,-4466,-15151,-17252,-5447,-9836,-1208,-3608,-9819,-11037,-3654,-14647,-5414,-8416,-3754,-8500,-8427,-2251,-8710,-2807,-2120,-3549,10762,3739,2519,3044,-3574,-6532,-2339,-6546,-6533,-11452,-8743,-3090,-5644,-2772,-8611,-6195,-10664,-8240,-14085,-9859,-14697,-5817,-4526,-2860,1518,1306,-7991,151,4420,5323,-3202,1141,-927,-8284,2417,-9049,-8237,-13733,-74,-3448,-1087,-6425,-10697,-3332,-12241,-13782,-5354,-7856,-12610,-12396,-9009,-7835,-6072,-2672,3263,-4109,-9323,-3252,-4716,-5673,1002,796,-3551,-5569,-3359,-4303,-5560,-11262,-11633,-14127,-14260,-5927,-12572,-7524,-12643,-18435,-13555,-7317,-5623,-492,-4957,-3763,2820,3379,-1689,-5186,-11043,479,-1639,-3689,4063,-2329,-8063,1022,-2387,-717,-6533,-14067,-8234,-8993,-13053,-14674,-3889,-11833,-15106,-2692,-2314,-2256,-3312,-7277,-2066,-4592,1888,-9810,473,-9455,-8637,-11284,-4430,-4458,1498,-1784,-6928,-1250,-4587,-5708,-3388,-9930,-8489,-9861,-6018,-12584,-5763,-1142,118,-6036,-5291,5280,-5969,-7817,-3173,-15218,-12627,-5283,4304,5565,-3528,6165,-924,-3957,2164,-9686,-4702,-10256,-13463,-15528,-3536,-14163,-13845,-2874,-9897,-9546,165,-8554,-1964,-3185,1763,-1815,-11488,-1596,-8672,53,274,4462,1256,-1529,4540,-6883,-3466,-1775,-12214,-7939,-5765,-15160,-16805,-14112,-14556,-16608,-11391,-7236,-6468,-5231,-8617,-2278,-7836,-9945,-4663,-3676,-6496,1070,9561,-2241,-3308,218,-1552,-7580,-2780,-2969,-15119,-3742,-1551,-9543,-15764,-16363,-17967,-13150,-7365,-4401,-5064,-9309,-11924,961,544,-3062,-2286,-7716,-7974,7046,8302,1810,223,-6681,-1509,-2932,-9593,-6088,-2063,-15087,-10819,-7835,-2763,-6077,-6596,-9575,-13190,-12860,1845,-13032,-448,-8377,-976,-5782,5179,-7785,-397,867,-1181,5268,-2571,305,-2716,-4774,-5802,-7907,-3215,-12088,-11671,-547,-13010,-12310,-8339,-10661,-5551,-12627,-5825,-11623,-8796,-8215,-7659,-10971,356,-5822,-3868,-2132,1609,-4691,-7312,1158,411,-13113,-7872,-13043,-14305,-10013,-11711,-14374,-5425,-12964,-7362,-13695,-10597,-16004,-8970,-12274,-4899,-14317,-3794,-10108,1570,-8512,-6378,507,-6526,-8180,-6945,2174,-1696,-12858,-2787,-2290,-7544,-7137,-5096,-6735,-2014,-15507,-5182,-8931,-9809,-9561,-6502,-17470,-15203,-14200,-14306,-6788,1896,166,136,1934,4446,-1638,1480,-7169,-2875,-3372,-9937,-12533,-3169,-2472,-1447,-9083,-6908,-12920,-3804,-2545,-5986,-17919,-11052,-11561,-2629,-10727,-8455,-6452,-8558,-1429,965,-3475,-11167,-667,-8979,-11579,-3615,-13431,-10669,-4439,-8558
};
layer_S #(18, 36, 15, 20, 784) L6(clk,reset,x,W,b,y,done);
endmodule